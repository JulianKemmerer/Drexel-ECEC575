# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2011, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on server08.nangate.com for user Giancarlo Franciscatto (gfr).
# Local time is now Thu, 6 Jan 2011, 18:10:28.
# Main process id is 3320.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO AON_BUF_X1
  CLASS core ;
  FOREIGN AON_BUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 1.33 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0378 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1586 LAYER metal1 ;
    ANTENNAGATEAREA 0.011 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.28 0.32 0.28 0.32 0.455 0.615 0.455 0.615 0.525 0.25 0.525  ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.04445 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1833 LAYER metal1 ;
    ANTENNADIFFAREA 0.0242 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.82 0.155 0.89 0.155 0.89 0.79 0.82 0.79  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.755 1.315 1.33 1.315 1.33 1.485 0.755 1.485 0 1.485  ;
    END
  END VDD
  PIN VDDBAK
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.92 0.595 0.92 0.595 0.735 0.73 0.735 0.73 0.92 0.755 0.92 0.94 0.92 0.94 1.12 0.755 1.12 0.385 1.12  ;
    END
  END VDDBAK
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 0.73 0.085 0.73 0.25 0.595 0.25 0.595 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.44 0.595 0.685 0.595 0.685 0.385 0.44 0.385 0.44 0.155 0.51 0.155 0.51 0.315 0.755 0.315 0.755 0.665 0.51 0.665 0.51 0.79 0.44 0.79  ;
  END
END AON_BUF_X1

END LIBRARY
#
# End of file
#
