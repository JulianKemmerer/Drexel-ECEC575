# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2011, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on server08.nangate.com for user Giancarlo Franciscatto (gfr).
# Local time is now Thu, 6 Jan 2011, 18:10:28.
# Main process id is 3320.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO LS_LH_X1
  CLASS core ;
  FOREIGN LS_LH_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 2.09 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0161 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0663 LAYER metal1 ;
    ANTENNAGATEAREA 0.01125 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.205 0.42 0.32 0.42 0.32 0.56 0.205 0.56  ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.06615 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2639 LAYER metal1 ;
    ANTENNADIFFAREA 0.0336 ;
    PORT
      LAYER metal1 ;
        POLYGON 1.96 0.19 2.03 0.19 2.03 1.135 1.96 1.135  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 1.37 1.315 1.37 1.085 1.44 1.085 1.44 1.315 1.77 1.315 1.77 1.125 1.84 1.125 1.84 1.315 1.89 1.315 2.09 1.315 2.09 1.485 1.89 1.485 0 1.485  ;
    END
  END VDD
  PIN VDDL
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.92 0.59 0.92 0.59 0.675 0.66 0.675 0.66 0.92 0.855 0.92 0.855 1.12 0.385 1.12  ;
    END
  END VDDL
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.09 -0.085 2.09 0.085 1.845 0.085 1.845 0.28 1.77 0.28 1.77 0.085 1.445 0.085 1.445 0.29 1.375 0.29 1.375 0.085 0.66 0.085 0.66 0.28 0.59 0.28 0.59 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.395 0.15 0.465 0.15 0.465 0.35 0.97 0.35 0.97 0.42 0.465 0.42 0.465 0.77 0.395 0.77  ;
        POLYGON 0.74 0.66 1.045 0.66 1.045 0.25 0.755 0.25 0.755 0.18 1.115 0.18 1.115 0.495 1.36 0.495 1.36 0.565 1.115 0.565 1.115 0.73 0.74 0.73  ;
        POLYGON 1.185 0.69 1.43 0.69 1.43 0.425 1.185 0.425 1.185 0.165 1.255 0.165 1.255 0.355 1.5 0.355 1.5 0.76 1.255 0.76 1.255 1.19 1.185 1.19  ;
        POLYGON 1.32 0.84 1.565 0.84 1.565 0.165 1.635 0.165 1.635 0.405 1.89 0.405 1.89 0.54 1.635 0.54 1.635 1.185 1.565 1.185 1.565 0.975 1.32 0.975  ;
  END
END LS_LH_X1

END LIBRARY
#
# End of file
#
