// Created by ihdl
module HEADER_X1 (SLEEP);
  input SLEEP;

endmodule
