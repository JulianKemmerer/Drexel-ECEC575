# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2010, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr).
# Local time is now Fri, 3 Dec 2010, 19:32:18.
# Main process id is 27821.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO SDFFR_X1
  CLASS core ;
  FOREIGN SDFFR_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 4.75 BY 1.4 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 ;
    PORT
      LAYER metal1 ;
        POLYGON 4.24 0.56 4.365 0.56 4.365 0.7 4.24 0.7  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0147 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0637 LAYER metal1 ;
    ANTENNAGATEAREA 0.03525 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.82 0.84 0.925 0.84 0.925 0.98 0.82 0.98  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0651 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2366 LAYER metal1 ;
    ANTENNAGATEAREA 0.05775 ;
    PORT
      LAYER metal1 ;
        POLYGON 4.105 0.565 4.175 0.565 4.175 0.77 4.43 0.77 4.43 0.56 4.53 0.56 4.53 0.84 4.105 0.84  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.017575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0728 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 ;
    PORT
      LAYER metal1 ;
        POLYGON 3.67 0.655 3.765 0.655 3.765 0.84 3.67 0.84  ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0405 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1053 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 ;
    PORT
      LAYER metal1 ;
        POLYGON 1.77 0.66 1.995 0.66 1.995 0.84 1.77 0.84  ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.06225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2353 LAYER metal1 ;
    ANTENNADIFFAREA 0.109725 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.435 0.185 0.51 0.185 0.51 1.015 0.435 1.015  ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.0616 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER metal1 ;
    ANTENNADIFFAREA 0.109725 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.185 0.13 0.185 0.13 1.065 0.06 1.065  ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.21 1.315 0.21 1.24 0.345 1.24 0.345 1.315 0.74 1.315 0.74 1.24 0.875 1.24 0.875 1.315 1.15 1.315 1.15 1.205 1.22 1.205 1.22 1.315 1.41 1.315 1.84 1.315 1.84 1.06 1.975 1.06 1.975 1.315 2.4 1.315 2.4 0.995 2.47 0.995 2.47 1.315 3.27 1.315 3.27 1.08 3.34 1.08 3.34 1.315 3.585 1.315 3.64 1.315 3.64 1.08 3.71 1.08 3.71 1.315 4.125 1.315 4.4 1.315 4.4 1.045 4.47 1.045 4.47 1.315 4.665 1.315 4.75 1.315 4.75 1.485 4.665 1.485 4.125 1.485 3.585 1.485 1.41 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 4.75 -0.085 4.75 0.085 4.47 0.085 4.47 0.32 4.4 0.32 4.4 0.085 3.71 0.085 3.71 0.32 3.64 0.32 3.64 0.085 3.18 0.085 3.18 0.32 3.11 0.32 3.11 0.085 2.34 0.085 2.34 0.425 2.27 0.425 2.27 0.085 1.845 0.085 1.845 0.285 1.71 0.285 1.71 0.085 0.84 0.085 0.84 0.32 0.77 0.32 0.77 0.085 0.31 0.085 0.31 0.46 0.24 0.46 0.24 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.195 0.525 0.265 0.525 0.265 1.08 0.585 1.08 0.585 0.185 0.655 0.185 0.655 0.39 1.075 0.39 1.075 0.635 1.005 0.635 1.005 0.46 0.655 0.46 0.655 1.24 0.585 1.24 0.585 1.15 0.195 1.15  ;
        POLYGON 0.935 1.045 1.41 1.045 1.41 1.115 0.935 1.115  ;
        POLYGON 1.21 0.905 1.56 0.905 1.56 1.04 1.49 1.04 1.49 0.975 1.14 0.975 1.14 0.775 0.72 0.775 0.72 0.525 0.79 0.525 0.79 0.705 1.14 0.705 1.14 0.215 1.46 0.215 1.46 0.285 1.21 0.285  ;
        POLYGON 1.35 0.765 1.695 0.765 1.695 0.905 2.065 0.905 2.065 0.655 2.26 0.655 2.26 0.79 2.135 0.79 2.135 1.065 2.065 1.065 2.065 0.975 1.695 0.975 1.695 1.25 1.545 1.25 1.545 1.18 1.625 1.18 1.625 0.835 1.28 0.835 1.28 0.35 1.93 0.35 1.93 0.185 2 0.185 2 0.42 1.35 0.42  ;
        POLYGON 2.22 0.855 2.335 0.855 2.335 0.56 1.5 0.56 1.5 0.7 1.43 0.7 1.43 0.49 2.09 0.49 2.09 0.185 2.16 0.185 2.16 0.49 2.405 0.49 2.405 0.17 2.92 0.17 2.92 0.835 2.85 0.835 2.85 0.24 2.475 0.24 2.475 0.56 2.405 0.56 2.405 0.925 2.29 0.925 2.29 1.13 2.22 1.13  ;
        POLYGON 2.69 0.305 2.76 0.305 2.76 1.015 2.995 1.015 2.995 0.81 3.45 0.81 3.45 0.88 3.065 0.88 3.065 1.085 2.69 1.085  ;
        POLYGON 2.54 0.505 2.61 0.505 2.61 1.18 3.135 1.18 3.135 0.945 3.515 0.945 3.515 0.725 2.985 0.725 2.985 0.385 3.265 0.385 3.265 0.185 3.335 0.185 3.335 0.455 3.055 0.455 3.055 0.655 3.585 0.655 3.585 1.015 3.52 1.015 3.52 1.2 3.45 1.2 3.45 1.015 3.205 1.015 3.205 1.25 2.54 1.25  ;
        POLYGON 3.9 1.04 4.125 1.04 4.125 1.11 3.83 1.11 3.83 0.59 3.12 0.59 3.12 0.52 3.83 0.52 3.83 0.22 4.125 0.22 4.125 0.29 3.9 0.29  ;
        POLYGON 3.965 0.715 4.035 0.715 4.035 0.905 4.595 0.905 4.595 0.485 4.1 0.485 4.1 0.415 4.595 0.415 4.595 0.185 4.665 0.185 4.665 1.22 4.595 1.22 4.595 0.975 3.965 0.975  ;
  END
END SDFFR_X1

END LIBRARY
#
# End of file
#
