# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2011, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on server08.nangate.com for user Giancarlo Franciscatto (gfr).
# Local time is now Thu, 6 Jan 2011, 18:10:28.
# Main process id is 3320.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO LS_LHEN_X2
  CLASS core ;
  FOREIGN LS_LHEN_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 2.66 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.03325 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1417 LAYER metal1 ;
    ANTENNAGATEAREA 0.011 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.47 0.565 0.47 0.565 0.54 0.32 0.54 0.32 0.7 0.25 0.7  ;
    END
  END A
  PIN ISOLN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0238 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0806 LAYER metal1 ;
    ANTENNAGATEAREA 0.02225 ;
    PORT
      LAYER metal1 ;
        POLYGON 1.86 0.7 2.03 0.7 2.03 0.84 1.86 0.84  ;
    END
  END ISOLN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.06825 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2717 LAYER metal1 ;
    ANTENNADIFFAREA 0.04725 ;
    PORT
      LAYER metal1 ;
        POLYGON 2.53 0.21 2.6 0.21 2.6 1.185 2.53 1.185  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.705 1.315 1.22 1.315 1.435 1.315 1.435 1.155 1.505 1.155 1.505 1.315 1.965 1.315 1.965 1.05 2.035 1.05 2.035 1.315 2.315 1.315 2.315 1.125 2.45 1.125 2.45 1.315 2.46 1.315 2.66 1.315 2.66 1.485 2.46 1.485 1.22 1.485 0.705 1.485 0 1.485  ;
    END
  END VDD
  PIN VDDL
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.415 0.92 0.55 0.92 0.55 0.74 0.685 0.74 0.685 0.92 0.705 0.92 0.83 0.92 0.83 1.12 0.705 1.12 0.415 1.12  ;
    END
  END VDDL
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.66 -0.085 2.66 0.085 2.45 0.085 2.45 0.225 2.315 0.225 2.315 0.085 1.88 0.085 1.88 0.34 1.81 0.34 1.81 0.085 0.98 0.085 0.98 0.335 0.91 0.335 0.91 0.085 0.605 0.085 0.605 0.27 0.535 0.27 0.535 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.395 0.605 0.635 0.605 0.635 0.405 0.345 0.405 0.345 0.15 0.415 0.15 0.415 0.335 0.705 0.335 0.705 0.675 0.465 0.675 0.465 0.795 0.395 0.795  ;
        POLYGON 0.695 0.17 0.845 0.17 0.845 0.54 1.15 0.54 1.15 0.365 1.22 0.365 1.22 0.61 0.845 0.61 0.845 0.795 0.775 0.795 0.775 0.24 0.695 0.24  ;
        POLYGON 1.245 0.77 1.285 0.77 1.285 0.21 1.355 0.21 1.355 0.77 1.575 0.77 1.575 0.84 1.315 0.84 1.315 1.23 1.245 1.23  ;
        POLYGON 1.385 0.92 1.645 0.92 1.645 0.585 1.44 0.585 1.44 0.21 1.51 0.21 1.51 0.515 2.325 0.515 2.325 0.585 1.715 0.585 1.715 1.23 1.645 1.23 1.645 1.055 1.385 1.055  ;
        POLYGON 2.155 0.835 2.39 0.835 2.39 0.44 1.97 0.44 1.97 0.17 2.04 0.17 2.04 0.37 2.46 0.37 2.46 0.905 2.225 0.905 2.225 1.185 2.155 1.185  ;
  END
END LS_LHEN_X2

END LIBRARY
#
# End of file
#
