# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2011, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on server08.nangate.com for user Giancarlo Franciscatto (gfr).
# Local time is now Thu, 6 Jan 2011, 18:10:28.
# Main process id is 3320.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO LS_LHEN_X1
  CLASS core ;
  FOREIGN LS_LHEN_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 2.66 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0308 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1326 LAYER metal1 ;
    ANTENNAGATEAREA 0.014 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.47 0.53 0.47 0.53 0.54 0.32 0.54 0.32 0.7 0.25 0.7  ;
    END
  END A
  PIN ISOLN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.026325 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0858 LAYER metal1 ;
    ANTENNAGATEAREA 0.0275 ;
    PORT
      LAYER metal1 ;
        POLYGON 1.895 0.645 2.03 0.645 2.03 0.84 1.895 0.84  ;
    END
  END ISOLN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.07725 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2873 LAYER metal1 ;
    ANTENNADIFFAREA 0.0336 ;
    PORT
      LAYER metal1 ;
        POLYGON 2.53 0.16 2.605 0.16 2.605 1.19 2.53 1.19  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.695 1.315 1.215 1.315 1.425 1.315 1.425 1.155 1.495 1.155 1.495 1.315 1.955 1.315 1.955 1.05 2.04 1.05 2.04 1.315 2.32 1.315 2.32 1.08 2.455 1.08 2.455 1.315 2.46 1.315 2.66 1.315 2.66 1.485 2.46 1.485 1.215 1.485 0.695 1.485 0 1.485  ;
    END
  END VDD
  PIN VDDL
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.41 0.92 0.55 0.92 0.55 0.74 0.685 0.74 0.685 0.92 0.695 0.92 0.83 0.92 0.83 1.12 0.695 1.12 0.41 1.12  ;
    END
  END VDDL
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.66 -0.085 2.66 0.085 2.42 0.085 2.42 0.295 2.35 0.295 2.35 0.085 1.875 0.085 1.875 0.32 1.805 0.32 1.805 0.085 0.975 0.085 0.975 0.32 0.905 0.32 0.905 0.085 0.62 0.085 0.62 0.27 0.55 0.27 0.55 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.4 0.605 0.625 0.605 0.625 0.405 0.365 0.405 0.365 0.15 0.435 0.15 0.435 0.335 0.695 0.335 0.695 0.675 0.47 0.675 0.47 0.74 0.4 0.74  ;
        POLYGON 0.705 0.165 0.84 0.165 0.84 0.44 1.145 0.44 1.145 0.325 1.215 0.325 1.215 0.51 0.84 0.51 0.84 0.74 0.77 0.74 0.77 0.235 0.705 0.235  ;
        POLYGON 1.245 0.775 1.28 0.775 1.28 0.185 1.35 0.185 1.35 0.775 1.565 0.775 1.565 0.845 1.315 0.845 1.315 1.23 1.245 1.23  ;
        POLYGON 1.38 0.92 1.64 0.92 1.64 0.575 1.435 0.575 1.435 0.185 1.505 0.185 1.505 0.505 2.325 0.505 2.325 0.575 1.71 0.575 1.71 1.23 1.64 1.23 1.64 1.055 1.38 1.055  ;
        POLYGON 2.16 0.935 2.39 0.935 2.39 0.435 1.975 0.435 1.975 0.16 2.045 0.16 2.045 0.365 2.46 0.365 2.46 1.005 2.23 1.005 2.23 1.19 2.16 1.19  ;
  END
END LS_LHEN_X1

END LIBRARY
#
# End of file
#
