# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2010, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr).
# Local time is now Fri, 3 Dec 2010, 19:32:18.
# Main process id is 27821.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO DFFRS_X1
  CLASS core ;
  FOREIGN DFFRS_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 4.56 BY 1.4 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.04845 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1157 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 ;
    PORT
      LAYER metal1 ;
        POLYGON 4.12 0.585 4.31 0.585 4.31 0.84 4.12 0.84  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0203 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0741 LAYER metal1 ;
    ANTENNAGATEAREA 0.03525 ;
    PORT
      LAYER metal1 ;
        POLYGON 1.2 0.7 1.345 0.7 1.345 0.84 1.2 0.84  ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0126 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0598 LAYER metal1 ;
    ANTENNAGATEAREA 0.0615 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.8 0.7 0.89 0.7 0.89 0.84 0.8 0.84  ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.031175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0936 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 ;
    PORT
      LAYER metal1 ;
        POLYGON 4.24 0.28 4.385 0.28 4.385 0.495 4.24 0.495  ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.03325 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1417 LAYER metal1 ;
    ANTENNADIFFAREA 0.109725 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.4 0.51 0.4 0.51 0.875 0.44 0.875  ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.0623 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2496 LAYER metal1 ;
    ANTENNADIFFAREA 0.109725 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.185 0.13 0.185 0.13 1.075 0.06 1.075  ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.215 1.315 0.215 1.1 0.35 1.1 0.35 1.315 0.56 1.315 0.56 1.095 0.695 1.095 0.695 1.315 0.88 1.315 0.965 1.315 0.965 1.065 1.035 1.065 1.035 1.315 1.345 1.315 1.345 0.925 1.415 0.925 1.415 1.315 1.655 1.315 1.655 0.99 1.79 0.99 1.79 1.315 1.945 1.315 2.415 1.315 2.415 0.89 2.55 0.89 2.55 1.315 2.795 1.315 2.795 0.835 2.93 0.835 2.93 1.315 3.325 1.315 3.325 1.03 3.46 1.03 3.46 1.315 3.615 1.315 4.055 1.315 4.255 1.315 4.255 0.915 4.325 0.915 4.325 1.315 4.52 1.315 4.56 1.315 4.56 1.485 4.52 1.485 4.055 1.485 3.615 1.485 1.945 1.485 0.88 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 4.56 -0.085 4.56 0.085 4.36 0.085 4.36 0.16 4.225 0.16 4.225 0.085 3.27 0.085 3.27 0.285 3.135 0.285 3.135 0.085 2.55 0.085 2.55 0.285 2.415 0.285 2.415 0.085 1.605 0.085 1.605 0.285 1.47 0.285 1.47 0.085 1.07 0.085 1.07 0.285 0.935 0.285 0.935 0.085 0.35 0.085 0.35 0.2 0.215 0.2 0.215 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.27 0.96 0.88 0.96 0.88 1.03 0.2 1.03 0.2 0.265 0.695 0.265 0.695 0.335 0.27 0.335  ;
        POLYGON 0.595 0.555 0.95 0.555 0.95 0.35 1.9 0.35 1.9 0.425 1.025 0.425 1.025 0.925 1.26 0.925 1.26 0.995 0.955 0.995 0.955 0.625 0.595 0.625  ;
        POLYGON 1.505 0.855 1.945 0.855 1.945 1.075 1.875 1.075 1.875 0.925 1.575 0.925 1.575 1.075 1.505 1.075  ;
        POLYGON 1.09 0.495 2.065 0.495 2.065 0.185 2.135 0.185 2.135 1.085 2.065 1.085 2.065 0.63 1.09 0.63  ;
        POLYGON 2.345 0.485 2.825 0.485 2.825 0.3 2.895 0.3 2.895 0.485 3.545 0.485 3.545 0.555 2.415 0.555 2.415 0.755 2.705 0.755 2.705 1.07 2.635 1.07 2.635 0.825 2.345 0.825  ;
        POLYGON 3.175 0.895 3.615 0.895 3.615 1.115 3.545 1.115 3.545 0.965 3.245 0.965 3.245 1.115 3.175 1.115  ;
        POLYGON 2.5 0.62 3.76 0.62 3.76 0.285 3.83 0.285 3.83 0.62 3.92 0.62 3.92 1.115 3.85 1.115 3.85 0.69 2.5 0.69  ;
        POLYGON 3.02 0.76 3.75 0.76 3.75 1.18 3.985 1.18 3.985 0.22 3.69 0.22 3.69 0.46 3.62 0.46 3.62 0.42 2.98 0.42 2.98 0.235 2.76 0.235 2.76 0.42 2.275 0.42 2.275 1.235 1.955 1.235 1.955 1.165 2.205 1.165 2.205 0.35 2.69 0.35 2.69 0.165 3.05 0.165 3.05 0.35 3.62 0.35 3.62 0.15 4.055 0.15 4.055 1.25 3.68 1.25 3.68 0.83 3.09 0.83 3.09 1.07 3.02 1.07  ;
        POLYGON 4.45 0.185 4.52 0.185 4.52 1.25 4.45 1.25  ;
  END
END DFFRS_X1

END LIBRARY
#
# End of file
#
