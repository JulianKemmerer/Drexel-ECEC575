# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2011, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on server08.nangate.com for user Giancarlo Franciscatto (gfr).
# Local time is now Thu, 6 Jan 2011, 18:10:28.
# Main process id is 3320.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO LS_LHEN_X4
  CLASS core ;
  FOREIGN LS_LHEN_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 2.66 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0329 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1404 LAYER metal1 ;
    ANTENNAGATEAREA 0.009 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.47 0.56 0.47 0.56 0.54 0.32 0.54 0.32 0.7 0.25 0.7  ;
    END
  END A
  PIN ISOLN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0231 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.0185 ;
    PORT
      LAYER metal1 ;
        POLYGON 1.865 0.7 2.03 0.7 2.03 0.84 1.865 0.84  ;
    END
  END ISOLN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.07175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2847 LAYER metal1 ;
    ANTENNADIFFAREA 0.0987 ;
    PORT
      LAYER metal1 ;
        POLYGON 2.53 0.18 2.6 0.18 2.6 1.205 2.53 1.205  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.695 1.315 1.21 1.315 1.395 1.315 1.395 1.155 1.53 1.155 1.53 1.315 1.96 1.315 1.96 1.1 2.03 1.1 2.03 1.315 2.34 1.315 2.34 1.1 2.41 1.1 2.41 1.315 2.46 1.315 2.66 1.315 2.66 1.485 2.46 1.485 1.21 1.485 0.695 1.485 0 1.485  ;
    END
  END VDD
  PIN VDDL
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.41 0.92 0.555 0.92 0.555 0.74 0.69 0.74 0.69 0.92 0.695 0.92 0.825 0.92 0.825 1.12 0.695 1.12 0.41 1.12  ;
    END
  END VDDL
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.66 -0.085 2.66 0.085 2.44 0.085 2.44 0.245 2.305 0.245 2.305 0.085 1.875 0.085 1.875 0.335 1.805 0.335 1.805 0.085 0.975 0.085 0.975 0.345 0.905 0.345 0.905 0.085 0.605 0.085 0.605 0.27 0.535 0.27 0.535 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.395 0.605 0.625 0.605 0.625 0.405 0.35 0.405 0.35 0.15 0.42 0.15 0.42 0.335 0.695 0.335 0.695 0.675 0.465 0.675 0.465 0.83 0.395 0.83  ;
        POLYGON 0.695 0.175 0.84 0.175 0.84 0.5 1.14 0.5 1.14 0.38 1.21 0.38 1.21 0.57 0.84 0.57 0.84 0.83 0.77 0.83 0.77 0.245 0.695 0.245  ;
        POLYGON 1.235 0.745 1.28 0.745 1.28 0.2 1.35 0.2 1.35 0.745 1.555 0.745 1.555 0.82 1.305 0.82 1.305 1.245 1.235 1.245  ;
        POLYGON 1.375 0.905 1.46 0.905 1.46 0.965 1.62 0.965 1.62 0.54 1.435 0.54 1.435 0.2 1.505 0.2 1.505 0.47 2.32 0.47 2.32 0.54 1.69 0.54 1.69 1.245 1.62 1.245 1.62 1.05 1.375 1.05  ;
        POLYGON 2.15 0.945 2.39 0.945 2.39 0.395 1.96 0.395 1.96 0.155 2.03 0.155 2.03 0.325 2.46 0.325 2.46 1.015 2.22 1.015 2.22 1.225 2.15 1.225  ;
  END
END LS_LHEN_X4

END LIBRARY
#
# End of file
#
