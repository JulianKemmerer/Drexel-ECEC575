# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2010, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr).
# Local time is now Fri, 3 Dec 2010, 19:32:18.
# Main process id is 27821.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO DFFS_X1
  CLASS core ;
  FOREIGN DFFS_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 3.8 BY 1.4 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0238 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0806 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.34 0.56 0.51 0.56 0.51 0.7 0.34 0.7  ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0231 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.03525 ;
    PORT
      LAYER metal1 ;
        POLYGON 2.625 0.7 2.79 0.7 2.79 0.84 2.625 0.84  ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.026275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1001 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 ;
    PORT
      LAYER metal1 ;
        POLYGON 1.705 0.59 1.84 0.59 1.84 0.84 1.77 0.84 1.77 0.725 1.705 0.725  ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.08155 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2964 LAYER metal1 ;
    ANTENNADIFFAREA 0.109725 ;
    PORT
      LAYER metal1 ;
        POLYGON 3.575 0.185 3.645 0.185 3.645 0.56 3.74 0.56 3.74 0.7 3.645 0.7 3.645 1.16 3.575 1.16  ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.0651 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2353 LAYER metal1 ;
    ANTENNADIFFAREA 0.109725 ;
    PORT
      LAYER metal1 ;
        POLYGON 3.195 0.185 3.265 0.185 3.265 0.56 3.36 0.56 3.36 0.7 3.265 0.7 3.265 0.925 3.195 0.925  ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.225 1.315 0.225 0.9 0.295 0.9 0.295 1.315 0.57 1.315 1.015 1.315 1.015 0.94 1.085 0.94 1.085 1.315 1.41 1.315 1.41 0.885 1.48 0.885 1.48 1.315 1.485 1.315 1.755 1.315 1.755 0.905 1.825 0.905 1.825 1.315 2.48 1.315 2.48 1.065 2.615 1.065 2.615 1.315 2.77 1.315 2.855 1.315 2.855 1.005 2.925 1.005 2.925 1.315 3.38 1.315 3.38 1.205 3.45 1.205 3.45 1.315 3.505 1.315 3.8 1.315 3.8 1.485 3.505 1.485 2.925 1.485 2.77 1.485 1.485 1.485 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 3.8 -0.085 3.8 0.085 3.455 0.085 3.455 0.46 3.385 0.46 3.385 0.085 2.805 0.085 2.805 0.34 2.67 0.34 2.67 0.085 1.82 0.085 1.82 0.375 1.75 0.375 1.75 0.085 1.11 0.085 1.11 0.32 1.04 0.32 1.04 0.085 0.295 0.085 0.295 0.32 0.225 0.32 0.225 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.04 0.185 0.11 0.185 0.11 0.765 0.57 0.765 0.57 0.835 0.11 0.835 0.11 1.16 0.04 1.16  ;
        POLYGON 0.59 0.975 0.795 0.975 0.795 0.615 0.77 0.615 0.77 0.355 0.59 0.355 0.59 0.285 0.84 0.285 0.84 0.545 1.35 0.545 1.35 0.685 1.28 0.685 1.28 0.615 0.865 0.615 0.865 1.045 0.59 1.045  ;
        POLYGON 0.94 0.685 1.01 0.685 1.01 0.75 1.415 0.75 1.415 0.285 1.485 0.285 1.485 0.82 1.29 0.82 1.29 1.09 1.22 1.09 1.22 0.82 0.94 0.82  ;
        POLYGON 0.175 0.42 0.445 0.42 0.445 0.15 0.975 0.15 0.975 0.385 1.28 0.385 1.28 0.15 1.64 0.15 1.64 0.44 1.97 0.44 1.97 0.15 2.32 0.15 2.32 0.22 2.04 0.22 2.04 0.665 2.095 0.665 2.095 0.8 1.97 0.8 1.97 0.51 1.64 0.51 1.64 0.815 1.67 0.815 1.67 1.09 1.57 1.09 1.57 0.22 1.35 0.22 1.35 0.455 0.905 0.455 0.905 0.22 0.515 0.22 0.515 0.42 0.705 0.42 0.705 0.72 0.73 0.72 0.73 0.855 0.635 0.855 0.635 0.49 0.245 0.49 0.245 0.685 0.175 0.685  ;
        POLYGON 2.33 0.93 2.77 0.93 2.77 1.15 2.7 1.15 2.7 1 2.4 1 2.4 1.15 2.33 1.15  ;
        POLYGON 2.105 1.045 2.17 1.045 2.17 0.36 2.105 0.36 2.105 0.29 2.24 0.29 2.24 0.56 2.925 0.56 2.925 0.63 2.24 0.63 2.24 1.115 2.105 1.115  ;
        POLYGON 2.375 0.42 2.905 0.42 2.905 0.185 2.975 0.185 2.975 0.42 3.08 0.42 3.08 0.995 3.435 0.995 3.435 0.525 3.505 0.525 3.505 1.065 3.01 1.065 3.01 0.49 2.375 0.49  ;
  END
END DFFS_X1

END LIBRARY
#
# End of file
#
