# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2011, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on server08.nangate.com for user Giancarlo Franciscatto (gfr).
# Local time is now Thu, 6 Jan 2011, 18:10:28.
# Main process id is 3320.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO LS_HL_X4
  CLASS core ;
  FOREIGN LS_HL_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0702 LAYER metal1 ;
    ANTENNAGATEAREA 0.02 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.19 0.42 0.19 0.56 0.06 0.56  ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.07065 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2275 LAYER metal1 ;
    ANTENNADIFFAREA 0.1008 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.425 0.15 0.515 0.15 0.515 0.935 0.425 0.935  ;
    END
  END Z
  PIN VDDL
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.225 1.315 0.225 0.815 0.295 0.815 0.295 1.315 0.355 1.315 0.605 1.315 0.605 0.815 0.675 0.815 0.675 1.315 0.76 1.315 0.76 1.485 0.355 1.485 0 1.485  ;
    END
  END VDDL
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.675 0.085 0.675 0.36 0.605 0.36 0.605 0.085 0.295 0.085 0.295 0.22 0.225 0.22 0.225 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.68 0.285 0.68 0.285 0.355 0.045 0.355 0.045 0.18 0.115 0.18 0.115 0.285 0.355 0.285 0.355 0.75 0.115 0.75 0.115 1.075 0.045 1.075  ;
  END
END LS_HL_X4

END LIBRARY
#
# End of file
#
