// Created by ihdl
module HEADER_X2 (SLEEP);
  input SLEEP;

endmodule
