# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2010, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr).
# Local time is now Fri, 3 Dec 2010, 19:32:18.
# Main process id is 27821.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO INV_X16
  CLASS core ;
  FOREIGN INV_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 3.23 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.357 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3442 LAYER metal1 ;
    ANTENNAGATEAREA 0.836 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.095 0.525 0.165 0.525 0.165 1.05 1.2 1.05 1.2 0.525 1.27 0.525 1.27 1.05 2 1.05 2 0.525 2.07 0.525 2.07 1.05 3.025 1.05 3.025 0.525 3.095 0.525 3.095 1.12 0.095 1.12  ;
    END
  END A
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.7672 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1788 LAYER metal1 ;
    ANTENNADIFFAREA 1.1704 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.18 0.305 0.18 0.305 0.28 0.605 0.28 0.605 0.16 0.675 0.16 0.675 0.28 0.985 0.28 0.985 0.15 1.055 0.15 1.055 0.28 1.365 0.28 1.365 0.15 1.435 0.15 1.435 0.28 1.745 0.28 1.745 0.15 1.815 0.15 1.815 0.28 2.125 0.28 2.125 0.15 2.195 0.15 2.195 0.28 2.505 0.28 2.505 0.15 2.575 0.15 2.575 0.28 2.885 0.28 2.885 0.15 2.955 0.15 2.955 0.985 2.885 0.985 2.885 0.42 2.575 0.42 2.575 0.985 2.505 0.985 2.505 0.42 2.205 0.42 2.205 0.985 2.135 0.985 2.135 0.42 1.815 0.42 1.815 0.985 1.745 0.985 1.745 0.42 1.435 0.42 1.435 0.985 1.365 0.985 1.365 0.42 1.055 0.42 1.055 0.985 0.985 0.985 0.985 0.42 0.675 0.42 0.675 0.985 0.605 0.985 0.605 0.42 0.305 0.42 0.305 0.985 0.235 0.985  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.205 0.11 1.205 0.11 1.315 0.415 1.315 0.415 1.205 0.485 1.205 0.485 1.315 0.795 1.315 0.795 1.205 0.865 1.205 0.865 1.315 1.175 1.315 1.175 1.205 1.245 1.205 1.245 1.315 1.555 1.315 1.555 1.205 1.625 1.205 1.625 1.315 1.935 1.315 1.935 1.205 2.005 1.205 2.005 1.315 2.315 1.315 2.315 1.205 2.385 1.205 2.385 1.315 2.695 1.315 2.695 1.205 2.765 1.205 2.765 1.315 3.075 1.315 3.075 1.205 3.145 1.205 3.145 1.315 3.23 1.315 3.23 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 3.23 -0.085 3.23 0.085 3.145 0.085 3.145 0.365 3.075 0.365 3.075 0.085 2.765 0.085 2.765 0.21 2.695 0.21 2.695 0.085 2.385 0.085 2.385 0.21 2.315 0.21 2.315 0.085 2.005 0.085 2.005 0.21 1.935 0.21 1.935 0.085 1.625 0.085 1.625 0.21 1.555 0.21 1.555 0.085 1.245 0.085 1.245 0.21 1.175 0.21 1.175 0.085 0.865 0.085 0.865 0.21 0.795 0.21 0.795 0.085 0.485 0.085 0.485 0.21 0.415 0.21 0.415 0.085 0.11 0.085 0.11 0.365 0.04 0.365 0.04 0.085 0 0.085  ;
    END
  END VSS
END INV_X16

END LIBRARY
#
# End of file
#
