# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2010, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr).
# Local time is now Fri, 3 Dec 2010, 19:32:18.
# Main process id is 27821.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO NAND4_X4
  CLASS core ;
  FOREIGN NAND4_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 3.42 BY 1.4 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.018375 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0728 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.405 0.525 0.51 0.525 0.51 0.7 0.405 0.7  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 ;
    PORT
      LAYER metal1 ;
        POLYGON 1.17 0.525 1.27 0.525 1.27 0.7 1.17 0.7  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.01225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0637 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 ;
    PORT
      LAYER metal1 ;
        POLYGON 2.15 0.525 2.22 0.525 2.22 0.7 2.15 0.7  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.01225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0637 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 ;
    PORT
      LAYER metal1 ;
        POLYGON 2.91 0.525 2.98 0.525 2.98 0.7 2.91 0.7  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.6363 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5548 LAYER metal1 ;
    ANTENNADIFFAREA 0.9604 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.09 0.84 0.685 0.84 0.685 0.355 0.225 0.355 0.225 0.285 0.755 0.285 0.755 0.84 2.425 0.84 3.34 0.84 3.34 1.155 3.27 1.155 3.27 0.98 2.96 0.98 2.96 1.155 2.89 1.155 2.89 0.98 2.58 0.98 2.58 1.155 2.51 1.155 2.51 0.98 2.425 0.98 2.2 0.98 2.2 1.155 2.13 1.155 2.13 0.98 1.75 0.98 1.75 1.155 1.68 1.155 1.68 0.98 1.29 0.98 1.29 1.155 1.22 1.155 1.22 0.98 0.91 0.98 0.91 1.155 0.84 1.155 0.84 0.98 0.53 0.98 0.53 1.155 0.46 1.155 0.46 0.98 0.16 0.98 0.16 1.155 0.09 1.155  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.24 1.315 0.24 1.095 0.375 1.095 0.375 1.315 0.62 1.315 0.62 1.095 0.755 1.095 0.755 1.315 1 1.315 1 1.095 1.135 1.095 1.135 1.315 1.38 1.315 1.38 1.095 1.515 1.095 1.515 1.315 1.91 1.315 1.91 1.095 2.045 1.095 2.045 1.315 2.29 1.315 2.29 1.095 2.425 1.095 2.425 1.315 2.67 1.315 2.67 1.095 2.805 1.095 2.805 1.315 3.05 1.315 3.05 1.095 3.185 1.095 3.185 1.315 3.34 1.315 3.42 1.315 3.42 1.485 3.34 1.485 2.425 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 3.42 -0.085 3.42 0.085 3.185 0.085 3.185 0.3 3.05 0.3 3.05 0.085 2.805 0.085 2.805 0.3 2.67 0.3 2.67 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.09 0.15 1.67 0.15 1.67 0.46 1.6 0.46 1.6 0.22 0.91 0.22 0.91 0.46 0.84 0.46 0.84 0.22 0.16 0.22 0.16 0.46 0.09 0.46  ;
        POLYGON 1.005 0.285 1.515 0.285 1.515 0.525 1.91 0.525 1.91 0.285 2.425 0.285 2.425 0.355 2.045 0.355 2.045 0.595 1.38 0.595 1.38 0.355 1.005 0.355  ;
        POLYGON 1.76 0.15 2.58 0.15 2.58 0.39 2.89 0.39 2.89 0.185 2.96 0.185 2.96 0.39 3.27 0.39 3.27 0.185 3.34 0.185 3.34 0.46 2.51 0.46 2.51 0.22 1.83 0.22 1.83 0.46 1.76 0.46  ;
  END
END NAND4_X4

END LIBRARY
#
# End of file
#
