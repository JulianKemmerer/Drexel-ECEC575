// Created by ihdl
module HEADER_X4 (SLEEP);
  input SLEEP;

endmodule
