# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2010, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr).
# Local time is now Fri, 3 Dec 2010, 19:32:18.
# Main process id is 27821.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO AOI21_X1
  CLASS core ;
  FOREIGN AOI21_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 0.76 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.575 0.525 0.7 0.525 0.7 0.7 0.575 0.7  ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.01925 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0741 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4 0.525 0.51 0.525 0.51 0.7 0.4 0.7  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0245 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0819 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.525 0.2 0.525 0.2 0.7 0.06 0.7  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.083925 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3185 LAYER metal1 ;
    ANTENNADIFFAREA 0.1463 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.265 0.355 0.44 0.355 0.44 0.15 0.525 0.15 0.525 0.425 0.335 0.425 0.335 1.115 0.265 1.115  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.525 1.315 0.645 1.315 0.645 0.905 0.715 0.905 0.715 1.315 0.76 1.315 0.76 1.485 0.525 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.715 0.085 0.715 0.355 0.645 0.355 0.645 0.085 0.15 0.085 0.15 0.425 0.08 0.425 0.08 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.085 0.905 0.155 0.905 0.155 1.18 0.455 1.18 0.455 0.905 0.525 0.905 0.525 1.25 0.085 1.25  ;
  END
END AOI21_X1

END LIBRARY
#
# End of file
#
