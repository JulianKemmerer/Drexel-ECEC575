# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2011, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on server08.nangate.com for user Giancarlo Franciscatto (gfr).
# Local time is now Thu, 6 Jan 2011, 18:10:28.
# Main process id is 3320.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO LS_HLEN_X4
  CLASS core ;
  FOREIGN LS_HLEN_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.02125 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0767 LAYER metal1 ;
    ANTENNAGATEAREA 0.0365 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.185 0.42 0.185 0.59 0.06 0.59  ;
    END
  END A
  PIN ISOLN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.02635 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0845 LAYER metal1 ;
    ANTENNAGATEAREA 0.0365 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.42 0.405 0.42 0.405 0.59 0.25 0.59  ;
    END
  END ISOLN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.0539 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2184 LAYER metal1 ;
    ANTENNADIFFAREA 0.1008 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.15 0.7 0.15 0.7 0.92 0.63 0.92  ;
    END
  END Z
  PIN VDDL
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.065 1.315 0.065 0.79 0.135 0.79 0.135 1.315 0.44 1.315 0.44 0.79 0.51 0.79 0.51 1.315 0.56 1.315 0.82 1.315 0.82 0.815 0.89 0.815 0.89 1.315 0.95 1.315 0.95 1.485 0.56 1.485 0 1.485  ;
    END
  END VDDL
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.89 0.085 0.89 0.34 0.82 0.34 0.82 0.085 0.51 0.085 0.51 0.2 0.44 0.2 0.44 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.26 0.655 0.49 0.655 0.49 0.355 0.035 0.355 0.035 0.285 0.56 0.285 0.56 0.725 0.33 0.725 0.33 0.93 0.26 0.93  ;
  END
END LS_HLEN_X4

END LIBRARY
#
# End of file
#
