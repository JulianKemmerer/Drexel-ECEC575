# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2010, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr).
# Local time is now Fri, 3 Dec 2010, 19:32:18.
# Main process id is 27821.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO AOI211_X4
  CLASS core ;
  FOREIGN AOI211_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 2.09 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.525 0.76 0.525 0.76 0.7 0.63 0.7  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.525 0.565 0.525 0.565 0.7 0.44 0.7  ;
    END
  END B
  PIN C1
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.525 0.185 0.525 0.185 0.7 0.06 0.7  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.525 0.375 0.525 0.375 0.7 0.25 0.7  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.1862 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6123 LAYER metal1 ;
    ANTENNADIFFAREA 0.2926 ;
    PORT
      LAYER metal1 ;
        POLYGON 1.375 0.15 1.445 0.15 1.445 0.56 1.75 0.56 1.75 0.15 1.82 0.15 1.82 1.175 1.75 1.175 1.75 0.7 1.445 0.7 1.445 1.175 1.375 1.175  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.485 1.315 0.795 1.315 0.795 0.9 0.865 0.9 0.865 1.315 0.93 1.315 1.175 1.315 1.175 0.9 1.245 0.9 1.245 1.315 1.31 1.315 1.555 1.315 1.555 0.9 1.625 0.9 1.625 1.315 1.935 1.315 1.935 0.9 2.005 0.9 2.005 1.315 2.09 1.315 2.09 1.485 1.31 1.485 0.93 1.485 0.485 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.09 -0.085 2.09 0.085 2.005 0.085 2.005 0.425 1.935 0.425 1.935 0.085 1.625 0.085 1.625 0.425 1.555 0.425 1.555 0.085 1.245 0.085 1.245 0.425 1.175 0.425 1.175 0.085 0.865 0.085 0.865 0.285 0.795 0.285 0.795 0.085 0.485 0.085 0.485 0.285 0.415 0.285 0.415 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.9 0.115 0.9 0.115 1.18 0.415 1.18 0.415 0.9 0.485 0.9 0.485 1.25 0.045 1.25  ;
        POLYGON 0.235 0.765 0.86 0.765 0.86 0.46 0.045 0.46 0.045 0.15 0.115 0.15 0.115 0.39 0.605 0.39 0.605 0.15 0.675 0.15 0.675 0.39 0.93 0.39 0.93 0.835 0.305 0.835 0.305 1.115 0.235 1.115  ;
        POLYGON 0.995 0.15 1.065 0.15 1.065 0.525 1.31 0.525 1.31 0.66 1.065 0.66 1.065 1.175 0.995 1.175  ;
  END
END AOI211_X4

END LIBRARY
#
# End of file
#
