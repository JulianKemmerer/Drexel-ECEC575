module add_unsigned_1245_GENERIC_REAL(A, B, Z);
// synthesis_equation add_unsigned
  input [52:0] A, B;
  output [52:0] Z;
  wire [52:0] A, B;
  wire [52:0] Z;
  wire n_161, n_166, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190;
  wire n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198;
  wire n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206;
  wire n_207, n_208, n_209, n_210, n_211, n_212, n_213, n_214;
  wire n_215, n_216, n_217, n_218, n_219, n_220, n_221, n_222;
  wire n_223, n_224, n_225, n_226, n_227, n_228, n_229, n_230;
  wire n_231, n_232, n_233, n_234, n_235, n_236, n_237, n_238;
  wire n_239, n_240, n_241, n_242, n_243, n_244, n_245, n_246;
  wire n_247, n_248, n_249, n_250, n_251, n_252, n_253, n_254;
  wire n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_262;
  wire n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270;
  wire n_271, n_272, n_273, n_274, n_275, n_276, n_277, n_278;
  wire n_279, n_280, n_281, n_282, n_283, n_284, n_285, n_286;
  wire n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_294;
  wire n_295, n_296, n_297, n_298, n_299, n_300, n_301, n_302;
  wire n_303, n_304, n_305, n_306, n_307, n_308, n_309, n_310;
  wire n_311, n_312, n_313, n_314, n_315, n_316, n_317, n_318;
  wire n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326;
  wire n_327, n_328, n_329, n_330, n_331, n_332, n_333, n_334;
  wire n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342;
  wire n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350;
  wire n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358;
  wire n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366;
  wire n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374;
  wire n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382;
  wire n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390;
  wire n_391, n_392, n_393, n_394, n_395, n_396, n_397, n_398;
  wire n_399, n_400, n_401, n_402, n_403, n_404, n_405, n_406;
  wire n_407, n_408, n_409, n_410, n_411, n_412, n_413, n_414;
  wire n_415, n_416, n_417, n_418, n_419, n_420, n_424, n_430;
  wire n_431;
  nand g1 (n_161, A[0], B[0]);
  xor g5 (Z[0], A[0], B[0]);
  nand g7 (n_166, A[1], B[1]);
  nand g10 (n_170, n_166, n_430, n_431);
  xor g11 (n_169, A[1], B[1]);
  nand g13 (n_171, A[2], B[2]);
  nand g14 (n_172, A[2], n_170);
  nand g15 (n_173, B[2], n_170);
  nand g16 (n_175, n_171, n_172, n_173);
  xor g17 (n_174, A[2], B[2]);
  xor g18 (Z[2], n_170, n_174);
  nand g19 (n_176, A[3], B[3]);
  nand g20 (n_177, A[3], n_175);
  nand g21 (n_178, B[3], n_175);
  nand g22 (n_180, n_176, n_177, n_178);
  xor g23 (n_179, A[3], B[3]);
  xor g24 (Z[3], n_175, n_179);
  nand g25 (n_181, A[4], B[4]);
  nand g26 (n_182, A[4], n_180);
  nand g27 (n_183, B[4], n_180);
  nand g28 (n_185, n_181, n_182, n_183);
  xor g29 (n_184, A[4], B[4]);
  xor g30 (Z[4], n_180, n_184);
  nand g31 (n_186, A[5], B[5]);
  nand g32 (n_187, A[5], n_185);
  nand g33 (n_188, B[5], n_185);
  nand g34 (n_190, n_186, n_187, n_188);
  xor g35 (n_189, A[5], B[5]);
  xor g36 (Z[5], n_185, n_189);
  nand g37 (n_191, A[6], B[6]);
  nand g38 (n_192, A[6], n_190);
  nand g39 (n_193, B[6], n_190);
  nand g40 (n_195, n_191, n_192, n_193);
  xor g41 (n_194, A[6], B[6]);
  xor g42 (Z[6], n_190, n_194);
  nand g43 (n_196, A[7], B[7]);
  nand g44 (n_197, A[7], n_195);
  nand g45 (n_198, B[7], n_195);
  nand g46 (n_200, n_196, n_197, n_198);
  xor g47 (n_199, A[7], B[7]);
  xor g48 (Z[7], n_195, n_199);
  nand g49 (n_201, A[8], B[8]);
  nand g50 (n_202, A[8], n_200);
  nand g51 (n_203, B[8], n_200);
  nand g52 (n_205, n_201, n_202, n_203);
  xor g53 (n_204, A[8], B[8]);
  xor g54 (Z[8], n_200, n_204);
  nand g55 (n_206, A[9], B[9]);
  nand g56 (n_207, A[9], n_205);
  nand g57 (n_208, B[9], n_205);
  nand g58 (n_210, n_206, n_207, n_208);
  xor g59 (n_209, A[9], B[9]);
  xor g60 (Z[9], n_205, n_209);
  nand g61 (n_211, A[10], B[10]);
  nand g62 (n_212, A[10], n_210);
  nand g63 (n_213, B[10], n_210);
  nand g64 (n_215, n_211, n_212, n_213);
  xor g65 (n_214, A[10], B[10]);
  xor g66 (Z[10], n_210, n_214);
  nand g67 (n_216, A[11], B[11]);
  nand g68 (n_217, A[11], n_215);
  nand g69 (n_218, B[11], n_215);
  nand g70 (n_220, n_216, n_217, n_218);
  xor g71 (n_219, A[11], B[11]);
  xor g72 (Z[11], n_215, n_219);
  nand g73 (n_221, A[12], B[12]);
  nand g74 (n_222, A[12], n_220);
  nand g75 (n_223, B[12], n_220);
  nand g76 (n_225, n_221, n_222, n_223);
  xor g77 (n_224, A[12], B[12]);
  xor g78 (Z[12], n_220, n_224);
  nand g79 (n_226, A[13], B[13]);
  nand g80 (n_227, A[13], n_225);
  nand g81 (n_228, B[13], n_225);
  nand g82 (n_230, n_226, n_227, n_228);
  xor g83 (n_229, A[13], B[13]);
  xor g84 (Z[13], n_225, n_229);
  nand g85 (n_231, A[14], B[14]);
  nand g86 (n_232, A[14], n_230);
  nand g87 (n_233, B[14], n_230);
  nand g88 (n_235, n_231, n_232, n_233);
  xor g89 (n_234, A[14], B[14]);
  xor g90 (Z[14], n_230, n_234);
  nand g91 (n_236, A[15], B[15]);
  nand g92 (n_237, A[15], n_235);
  nand g93 (n_238, B[15], n_235);
  nand g94 (n_240, n_236, n_237, n_238);
  xor g95 (n_239, A[15], B[15]);
  xor g96 (Z[15], n_235, n_239);
  nand g97 (n_241, A[16], B[16]);
  nand g98 (n_242, A[16], n_240);
  nand g99 (n_243, B[16], n_240);
  nand g100 (n_245, n_241, n_242, n_243);
  xor g101 (n_244, A[16], B[16]);
  xor g102 (Z[16], n_240, n_244);
  nand g103 (n_246, A[17], B[17]);
  nand g104 (n_247, A[17], n_245);
  nand g105 (n_248, B[17], n_245);
  nand g106 (n_250, n_246, n_247, n_248);
  xor g107 (n_249, A[17], B[17]);
  xor g108 (Z[17], n_245, n_249);
  nand g109 (n_251, A[18], B[18]);
  nand g110 (n_252, A[18], n_250);
  nand g111 (n_253, B[18], n_250);
  nand g112 (n_255, n_251, n_252, n_253);
  xor g113 (n_254, A[18], B[18]);
  xor g114 (Z[18], n_250, n_254);
  nand g115 (n_256, A[19], B[19]);
  nand g116 (n_257, A[19], n_255);
  nand g117 (n_258, B[19], n_255);
  nand g118 (n_260, n_256, n_257, n_258);
  xor g119 (n_259, A[19], B[19]);
  xor g120 (Z[19], n_255, n_259);
  nand g121 (n_261, A[20], B[20]);
  nand g122 (n_262, A[20], n_260);
  nand g123 (n_263, B[20], n_260);
  nand g124 (n_265, n_261, n_262, n_263);
  xor g125 (n_264, A[20], B[20]);
  xor g126 (Z[20], n_260, n_264);
  nand g127 (n_266, A[21], B[21]);
  nand g128 (n_267, A[21], n_265);
  nand g129 (n_268, B[21], n_265);
  nand g130 (n_270, n_266, n_267, n_268);
  xor g131 (n_269, A[21], B[21]);
  xor g132 (Z[21], n_265, n_269);
  nand g133 (n_271, A[22], B[22]);
  nand g134 (n_272, A[22], n_270);
  nand g135 (n_273, B[22], n_270);
  nand g136 (n_275, n_271, n_272, n_273);
  xor g137 (n_274, A[22], B[22]);
  xor g138 (Z[22], n_270, n_274);
  nand g139 (n_276, A[23], B[23]);
  nand g140 (n_277, A[23], n_275);
  nand g141 (n_278, B[23], n_275);
  nand g142 (n_280, n_276, n_277, n_278);
  xor g143 (n_279, A[23], B[23]);
  xor g144 (Z[23], n_275, n_279);
  nand g145 (n_281, A[24], B[24]);
  nand g146 (n_282, A[24], n_280);
  nand g147 (n_283, B[24], n_280);
  nand g148 (n_285, n_281, n_282, n_283);
  xor g149 (n_284, A[24], B[24]);
  xor g150 (Z[24], n_280, n_284);
  nand g151 (n_286, A[25], B[25]);
  nand g152 (n_287, A[25], n_285);
  nand g153 (n_288, B[25], n_285);
  nand g154 (n_290, n_286, n_287, n_288);
  xor g155 (n_289, A[25], B[25]);
  xor g156 (Z[25], n_285, n_289);
  nand g157 (n_291, A[26], B[26]);
  nand g158 (n_292, A[26], n_290);
  nand g159 (n_293, B[26], n_290);
  nand g160 (n_295, n_291, n_292, n_293);
  xor g161 (n_294, A[26], B[26]);
  xor g162 (Z[26], n_290, n_294);
  nand g163 (n_296, A[27], B[27]);
  nand g164 (n_297, A[27], n_295);
  nand g165 (n_298, B[27], n_295);
  nand g166 (n_300, n_296, n_297, n_298);
  xor g167 (n_299, A[27], B[27]);
  xor g168 (Z[27], n_295, n_299);
  nand g169 (n_301, A[28], B[28]);
  nand g170 (n_302, A[28], n_300);
  nand g171 (n_303, B[28], n_300);
  nand g172 (n_305, n_301, n_302, n_303);
  xor g173 (n_304, A[28], B[28]);
  xor g174 (Z[28], n_300, n_304);
  nand g175 (n_306, A[29], B[29]);
  nand g176 (n_307, A[29], n_305);
  nand g177 (n_308, B[29], n_305);
  nand g178 (n_310, n_306, n_307, n_308);
  xor g179 (n_309, A[29], B[29]);
  xor g180 (Z[29], n_305, n_309);
  nand g181 (n_311, A[30], B[30]);
  nand g182 (n_312, A[30], n_310);
  nand g183 (n_313, B[30], n_310);
  nand g184 (n_315, n_311, n_312, n_313);
  xor g185 (n_314, A[30], B[30]);
  xor g186 (Z[30], n_310, n_314);
  nand g187 (n_316, A[31], B[31]);
  nand g188 (n_317, A[31], n_315);
  nand g189 (n_318, B[31], n_315);
  nand g190 (n_320, n_316, n_317, n_318);
  xor g191 (n_319, A[31], B[31]);
  xor g192 (Z[31], n_315, n_319);
  nand g193 (n_321, A[32], B[32]);
  nand g194 (n_322, A[32], n_320);
  nand g195 (n_323, B[32], n_320);
  nand g196 (n_325, n_321, n_322, n_323);
  xor g197 (n_324, A[32], B[32]);
  xor g198 (Z[32], n_320, n_324);
  nand g199 (n_326, A[33], B[33]);
  nand g200 (n_327, A[33], n_325);
  nand g201 (n_328, B[33], n_325);
  nand g202 (n_330, n_326, n_327, n_328);
  xor g203 (n_329, A[33], B[33]);
  xor g204 (Z[33], n_325, n_329);
  nand g205 (n_331, A[34], B[34]);
  nand g206 (n_332, A[34], n_330);
  nand g207 (n_333, B[34], n_330);
  nand g208 (n_335, n_331, n_332, n_333);
  xor g209 (n_334, A[34], B[34]);
  xor g210 (Z[34], n_330, n_334);
  nand g211 (n_336, A[35], B[35]);
  nand g212 (n_337, A[35], n_335);
  nand g213 (n_338, B[35], n_335);
  nand g214 (n_340, n_336, n_337, n_338);
  xor g215 (n_339, A[35], B[35]);
  xor g216 (Z[35], n_335, n_339);
  nand g217 (n_341, A[36], B[36]);
  nand g218 (n_342, A[36], n_340);
  nand g219 (n_343, B[36], n_340);
  nand g220 (n_345, n_341, n_342, n_343);
  xor g221 (n_344, A[36], B[36]);
  xor g222 (Z[36], n_340, n_344);
  nand g223 (n_346, A[37], B[37]);
  nand g224 (n_347, A[37], n_345);
  nand g225 (n_348, B[37], n_345);
  nand g226 (n_350, n_346, n_347, n_348);
  xor g227 (n_349, A[37], B[37]);
  xor g228 (Z[37], n_345, n_349);
  nand g229 (n_351, A[38], B[38]);
  nand g230 (n_352, A[38], n_350);
  nand g231 (n_353, B[38], n_350);
  nand g232 (n_355, n_351, n_352, n_353);
  xor g233 (n_354, A[38], B[38]);
  xor g234 (Z[38], n_350, n_354);
  nand g235 (n_356, A[39], B[39]);
  nand g236 (n_357, A[39], n_355);
  nand g237 (n_358, B[39], n_355);
  nand g238 (n_360, n_356, n_357, n_358);
  xor g239 (n_359, A[39], B[39]);
  xor g240 (Z[39], n_355, n_359);
  nand g241 (n_361, A[40], B[40]);
  nand g242 (n_362, A[40], n_360);
  nand g243 (n_363, B[40], n_360);
  nand g244 (n_365, n_361, n_362, n_363);
  xor g245 (n_364, A[40], B[40]);
  xor g246 (Z[40], n_360, n_364);
  nand g247 (n_366, A[41], B[41]);
  nand g248 (n_367, A[41], n_365);
  nand g249 (n_368, B[41], n_365);
  nand g250 (n_370, n_366, n_367, n_368);
  xor g251 (n_369, A[41], B[41]);
  xor g252 (Z[41], n_365, n_369);
  nand g253 (n_371, A[42], B[42]);
  nand g254 (n_372, A[42], n_370);
  nand g255 (n_373, B[42], n_370);
  nand g256 (n_375, n_371, n_372, n_373);
  xor g257 (n_374, A[42], B[42]);
  xor g258 (Z[42], n_370, n_374);
  nand g259 (n_376, A[43], B[43]);
  nand g260 (n_377, A[43], n_375);
  nand g261 (n_378, B[43], n_375);
  nand g262 (n_380, n_376, n_377, n_378);
  xor g263 (n_379, A[43], B[43]);
  xor g264 (Z[43], n_375, n_379);
  nand g265 (n_381, A[44], B[44]);
  nand g266 (n_382, A[44], n_380);
  nand g267 (n_383, B[44], n_380);
  nand g268 (n_385, n_381, n_382, n_383);
  xor g269 (n_384, A[44], B[44]);
  xor g270 (Z[44], n_380, n_384);
  nand g271 (n_386, A[45], B[45]);
  nand g272 (n_387, A[45], n_385);
  nand g273 (n_388, B[45], n_385);
  nand g274 (n_390, n_386, n_387, n_388);
  xor g275 (n_389, A[45], B[45]);
  xor g276 (Z[45], n_385, n_389);
  nand g277 (n_391, A[46], B[46]);
  nand g278 (n_392, A[46], n_390);
  nand g279 (n_393, B[46], n_390);
  nand g280 (n_395, n_391, n_392, n_393);
  xor g281 (n_394, A[46], B[46]);
  xor g282 (Z[46], n_390, n_394);
  nand g283 (n_396, A[47], B[47]);
  nand g284 (n_397, A[47], n_395);
  nand g285 (n_398, B[47], n_395);
  nand g286 (n_400, n_396, n_397, n_398);
  xor g287 (n_399, A[47], B[47]);
  xor g288 (Z[47], n_395, n_399);
  nand g289 (n_401, A[48], B[48]);
  nand g290 (n_402, A[48], n_400);
  nand g291 (n_403, B[48], n_400);
  nand g292 (n_405, n_401, n_402, n_403);
  xor g293 (n_404, A[48], B[48]);
  xor g294 (Z[48], n_400, n_404);
  nand g295 (n_406, A[49], B[49]);
  nand g296 (n_407, A[49], n_405);
  nand g297 (n_408, B[49], n_405);
  nand g298 (n_410, n_406, n_407, n_408);
  xor g299 (n_409, A[49], B[49]);
  xor g300 (Z[49], n_405, n_409);
  nand g301 (n_411, A[50], B[50]);
  nand g302 (n_412, A[50], n_410);
  nand g303 (n_413, B[50], n_410);
  nand g304 (n_415, n_411, n_412, n_413);
  xor g305 (n_414, A[50], B[50]);
  xor g306 (Z[50], n_410, n_414);
  nand g307 (n_416, A[51], B[51]);
  nand g308 (n_417, A[51], n_415);
  nand g309 (n_418, B[51], n_415);
  nand g310 (n_420, n_416, n_417, n_418);
  xor g311 (n_419, A[51], B[51]);
  xor g312 (Z[51], n_415, n_419);
  xor g317 (n_424, A[52], B[52]);
  xor g318 (Z[52], n_420, n_424);
  or g320 (n_430, wc, n_161);
  not gc (wc, A[1]);
  or g321 (n_431, wc0, n_161);
  not gc0 (wc0, B[1]);
  xnor g322 (Z[1], n_161, n_169);
endmodule

module add_unsigned_1245_GENERIC(A, B, Z);
  input [52:0] A, B;
  output [52:0] Z;
  wire [52:0] A, B;
  wire [52:0] Z;
  add_unsigned_1245_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_unsigned_2994_GENERIC_REAL(A, B, Z);
// synthesis_equation add_unsigned
  input [32:0] A, B;
  output [32:0] Z;
  wire [32:0] A, B;
  wire [32:0] Z;
  wire n_101, n_106, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_264, n_270, n_271;
  nand g1 (n_101, A[0], B[0]);
  xor g5 (Z[0], A[0], B[0]);
  nand g7 (n_106, A[1], B[1]);
  nand g10 (n_110, n_106, n_270, n_271);
  xor g11 (n_109, A[1], B[1]);
  nand g13 (n_111, A[2], B[2]);
  nand g14 (n_112, A[2], n_110);
  nand g15 (n_113, B[2], n_110);
  nand g16 (n_115, n_111, n_112, n_113);
  xor g17 (n_114, A[2], B[2]);
  xor g18 (Z[2], n_110, n_114);
  nand g19 (n_116, A[3], B[3]);
  nand g20 (n_117, A[3], n_115);
  nand g21 (n_118, B[3], n_115);
  nand g22 (n_120, n_116, n_117, n_118);
  xor g23 (n_119, A[3], B[3]);
  xor g24 (Z[3], n_115, n_119);
  nand g25 (n_121, A[4], B[4]);
  nand g26 (n_122, A[4], n_120);
  nand g27 (n_123, B[4], n_120);
  nand g28 (n_125, n_121, n_122, n_123);
  xor g29 (n_124, A[4], B[4]);
  xor g30 (Z[4], n_120, n_124);
  nand g31 (n_126, A[5], B[5]);
  nand g32 (n_127, A[5], n_125);
  nand g33 (n_128, B[5], n_125);
  nand g34 (n_130, n_126, n_127, n_128);
  xor g35 (n_129, A[5], B[5]);
  xor g36 (Z[5], n_125, n_129);
  nand g37 (n_131, A[6], B[6]);
  nand g38 (n_132, A[6], n_130);
  nand g39 (n_133, B[6], n_130);
  nand g40 (n_135, n_131, n_132, n_133);
  xor g41 (n_134, A[6], B[6]);
  xor g42 (Z[6], n_130, n_134);
  nand g43 (n_136, A[7], B[7]);
  nand g44 (n_137, A[7], n_135);
  nand g45 (n_138, B[7], n_135);
  nand g46 (n_140, n_136, n_137, n_138);
  xor g47 (n_139, A[7], B[7]);
  xor g48 (Z[7], n_135, n_139);
  nand g49 (n_141, A[8], B[8]);
  nand g50 (n_142, A[8], n_140);
  nand g51 (n_143, B[8], n_140);
  nand g52 (n_145, n_141, n_142, n_143);
  xor g53 (n_144, A[8], B[8]);
  xor g54 (Z[8], n_140, n_144);
  nand g55 (n_146, A[9], B[9]);
  nand g56 (n_147, A[9], n_145);
  nand g57 (n_148, B[9], n_145);
  nand g58 (n_150, n_146, n_147, n_148);
  xor g59 (n_149, A[9], B[9]);
  xor g60 (Z[9], n_145, n_149);
  nand g61 (n_151, A[10], B[10]);
  nand g62 (n_152, A[10], n_150);
  nand g63 (n_153, B[10], n_150);
  nand g64 (n_155, n_151, n_152, n_153);
  xor g65 (n_154, A[10], B[10]);
  xor g66 (Z[10], n_150, n_154);
  nand g67 (n_156, A[11], B[11]);
  nand g68 (n_157, A[11], n_155);
  nand g69 (n_158, B[11], n_155);
  nand g70 (n_160, n_156, n_157, n_158);
  xor g71 (n_159, A[11], B[11]);
  xor g72 (Z[11], n_155, n_159);
  nand g73 (n_161, A[12], B[12]);
  nand g74 (n_162, A[12], n_160);
  nand g75 (n_163, B[12], n_160);
  nand g76 (n_165, n_161, n_162, n_163);
  xor g77 (n_164, A[12], B[12]);
  xor g78 (Z[12], n_160, n_164);
  nand g79 (n_166, A[13], B[13]);
  nand g80 (n_167, A[13], n_165);
  nand g81 (n_168, B[13], n_165);
  nand g82 (n_170, n_166, n_167, n_168);
  xor g83 (n_169, A[13], B[13]);
  xor g84 (Z[13], n_165, n_169);
  nand g85 (n_171, A[14], B[14]);
  nand g86 (n_172, A[14], n_170);
  nand g87 (n_173, B[14], n_170);
  nand g88 (n_175, n_171, n_172, n_173);
  xor g89 (n_174, A[14], B[14]);
  xor g90 (Z[14], n_170, n_174);
  nand g91 (n_176, A[15], B[15]);
  nand g92 (n_177, A[15], n_175);
  nand g93 (n_178, B[15], n_175);
  nand g94 (n_180, n_176, n_177, n_178);
  xor g95 (n_179, A[15], B[15]);
  xor g96 (Z[15], n_175, n_179);
  nand g97 (n_181, A[16], B[16]);
  nand g98 (n_182, A[16], n_180);
  nand g99 (n_183, B[16], n_180);
  nand g100 (n_185, n_181, n_182, n_183);
  xor g101 (n_184, A[16], B[16]);
  xor g102 (Z[16], n_180, n_184);
  nand g103 (n_186, A[17], B[17]);
  nand g104 (n_187, A[17], n_185);
  nand g105 (n_188, B[17], n_185);
  nand g106 (n_190, n_186, n_187, n_188);
  xor g107 (n_189, A[17], B[17]);
  xor g108 (Z[17], n_185, n_189);
  nand g109 (n_191, A[18], B[18]);
  nand g110 (n_192, A[18], n_190);
  nand g111 (n_193, B[18], n_190);
  nand g112 (n_195, n_191, n_192, n_193);
  xor g113 (n_194, A[18], B[18]);
  xor g114 (Z[18], n_190, n_194);
  nand g115 (n_196, A[19], B[19]);
  nand g116 (n_197, A[19], n_195);
  nand g117 (n_198, B[19], n_195);
  nand g118 (n_200, n_196, n_197, n_198);
  xor g119 (n_199, A[19], B[19]);
  xor g120 (Z[19], n_195, n_199);
  nand g121 (n_201, A[20], B[20]);
  nand g122 (n_202, A[20], n_200);
  nand g123 (n_203, B[20], n_200);
  nand g124 (n_205, n_201, n_202, n_203);
  xor g125 (n_204, A[20], B[20]);
  xor g126 (Z[20], n_200, n_204);
  nand g127 (n_206, A[21], B[21]);
  nand g128 (n_207, A[21], n_205);
  nand g129 (n_208, B[21], n_205);
  nand g130 (n_210, n_206, n_207, n_208);
  xor g131 (n_209, A[21], B[21]);
  xor g132 (Z[21], n_205, n_209);
  nand g133 (n_211, A[22], B[22]);
  nand g134 (n_212, A[22], n_210);
  nand g135 (n_213, B[22], n_210);
  nand g136 (n_215, n_211, n_212, n_213);
  xor g137 (n_214, A[22], B[22]);
  xor g138 (Z[22], n_210, n_214);
  nand g139 (n_216, A[23], B[23]);
  nand g140 (n_217, A[23], n_215);
  nand g141 (n_218, B[23], n_215);
  nand g142 (n_220, n_216, n_217, n_218);
  xor g143 (n_219, A[23], B[23]);
  xor g144 (Z[23], n_215, n_219);
  nand g145 (n_221, A[24], B[24]);
  nand g146 (n_222, A[24], n_220);
  nand g147 (n_223, B[24], n_220);
  nand g148 (n_225, n_221, n_222, n_223);
  xor g149 (n_224, A[24], B[24]);
  xor g150 (Z[24], n_220, n_224);
  nand g151 (n_226, A[25], B[25]);
  nand g152 (n_227, A[25], n_225);
  nand g153 (n_228, B[25], n_225);
  nand g154 (n_230, n_226, n_227, n_228);
  xor g155 (n_229, A[25], B[25]);
  xor g156 (Z[25], n_225, n_229);
  nand g157 (n_231, A[26], B[26]);
  nand g158 (n_232, A[26], n_230);
  nand g159 (n_233, B[26], n_230);
  nand g160 (n_235, n_231, n_232, n_233);
  xor g161 (n_234, A[26], B[26]);
  xor g162 (Z[26], n_230, n_234);
  nand g163 (n_236, A[27], B[27]);
  nand g164 (n_237, A[27], n_235);
  nand g165 (n_238, B[27], n_235);
  nand g166 (n_240, n_236, n_237, n_238);
  xor g167 (n_239, A[27], B[27]);
  xor g168 (Z[27], n_235, n_239);
  nand g169 (n_241, A[28], B[28]);
  nand g170 (n_242, A[28], n_240);
  nand g171 (n_243, B[28], n_240);
  nand g172 (n_245, n_241, n_242, n_243);
  xor g173 (n_244, A[28], B[28]);
  xor g174 (Z[28], n_240, n_244);
  nand g175 (n_246, A[29], B[29]);
  nand g176 (n_247, A[29], n_245);
  nand g177 (n_248, B[29], n_245);
  nand g178 (n_250, n_246, n_247, n_248);
  xor g179 (n_249, A[29], B[29]);
  xor g180 (Z[29], n_245, n_249);
  nand g181 (n_251, A[30], B[30]);
  nand g182 (n_252, A[30], n_250);
  nand g183 (n_253, B[30], n_250);
  nand g184 (n_255, n_251, n_252, n_253);
  xor g185 (n_254, A[30], B[30]);
  xor g186 (Z[30], n_250, n_254);
  nand g187 (n_256, A[31], B[31]);
  nand g188 (n_257, A[31], n_255);
  nand g189 (n_258, B[31], n_255);
  nand g190 (n_260, n_256, n_257, n_258);
  xor g191 (n_259, A[31], B[31]);
  xor g192 (Z[31], n_255, n_259);
  xor g197 (n_264, A[32], B[32]);
  xor g198 (Z[32], n_260, n_264);
  or g200 (n_270, wc, n_101);
  not gc (wc, A[1]);
  or g201 (n_271, wc0, n_101);
  not gc0 (wc0, B[1]);
  xnor g202 (Z[1], n_101, n_109);
endmodule

module add_unsigned_2994_GENERIC(A, B, Z);
  input [32:0] A, B;
  output [32:0] Z;
  wire [32:0] A, B;
  wire [32:0] Z;
  add_unsigned_2994_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_unsigned_carry_2513_GENERIC_REAL(A, B, CI, Z);
// synthesis_equation add_unsigned_carry
  input [63:0] A, B;
  input CI;
  output [63:0] Z;
  wire [63:0] A, B;
  wire CI;
  wire [63:0] Z;
  wire n_194, n_195, n_196, n_197, n_198, n_200, n_202, n_203;
  wire n_204, n_205, n_207, n_208, n_209, n_210, n_211, n_213;
  wire n_214, n_215, n_216, n_217, n_219, n_220, n_221, n_222;
  wire n_223, n_225, n_226, n_227, n_228, n_229, n_231, n_232;
  wire n_233, n_234, n_235, n_237, n_238, n_239, n_240, n_241;
  wire n_243, n_244, n_245, n_246, n_247, n_249, n_250, n_251;
  wire n_252, n_253, n_255, n_256, n_257, n_258, n_259, n_261;
  wire n_262, n_263, n_264, n_265, n_267, n_268, n_269, n_270;
  wire n_271, n_273, n_274, n_275, n_276, n_277, n_279, n_280;
  wire n_281, n_282, n_283, n_285, n_286, n_287, n_288, n_289;
  wire n_291, n_292, n_293, n_294, n_295, n_297, n_298, n_299;
  wire n_300, n_301, n_303, n_304, n_305, n_306, n_307, n_309;
  wire n_310, n_311, n_312, n_313, n_315, n_316, n_317, n_318;
  wire n_319, n_321, n_322, n_323, n_324, n_325, n_327, n_328;
  wire n_329, n_330, n_331, n_333, n_334, n_335, n_336, n_337;
  wire n_339, n_340, n_341, n_342, n_343, n_345, n_346, n_347;
  wire n_348, n_349, n_351, n_352, n_353, n_354, n_355, n_357;
  wire n_358, n_359, n_360, n_361, n_363, n_364, n_365, n_366;
  wire n_367, n_369, n_370, n_371, n_372, n_373, n_375, n_376;
  wire n_377, n_378, n_379, n_381, n_382, n_383, n_384, n_387;
  wire n_388, n_389, n_391, n_392, n_393, n_398, n_399, n_400;
  wire n_405, n_406, n_407, n_412, n_413, n_414, n_419, n_420;
  wire n_421, n_426, n_427, n_428, n_433, n_434, n_435, n_440;
  wire n_441, n_442, n_447, n_448, n_449, n_454, n_455, n_456;
  wire n_461, n_462, n_463, n_468, n_469, n_470, n_475, n_476;
  wire n_477, n_482, n_483, n_484, n_489, n_496, n_497, n_498;
  wire n_502, n_503, n_505, n_507, n_508, n_509, n_511, n_513;
  wire n_514, n_515, n_517, n_519, n_520, n_521, n_523, n_525;
  wire n_526, n_527, n_529, n_531, n_532, n_533, n_535, n_537;
  wire n_543, n_544, n_545, n_547, n_548, n_549, n_554, n_555;
  wire n_556, n_561, n_568, n_569, n_570, n_579, n_581, n_586;
  wire n_587, n_588, n_589, n_594, n_599, n_604, n_607, n_608;
  wire n_609, n_610, n_611, n_612, n_613, n_614, n_615, n_616;
  wire n_617, n_618, n_619, n_620, n_621, n_622, n_623, n_624;
  wire n_625, n_626, n_627, n_628, n_633, n_638, n_643, n_648;
  wire n_653, n_658, n_663, n_668, n_673, n_678, n_683, n_688;
  wire n_693, n_698, n_703, n_709, n_713, n_717, n_721, n_725;
  wire n_729, n_733, n_737, n_741, n_745, n_749, n_753, n_757;
  wire n_761, n_765, n_769, n_773, n_777, n_781, n_785, n_789;
  wire n_793, n_797, n_801, n_805, n_809, n_813, n_817, n_821;
  wire n_825, n_829, n_831, n_837, n_838, n_839, n_840, n_841;
  wire n_842, n_843, n_844, n_845, n_846, n_847, n_848, n_849;
  wire n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857;
  wire n_858, n_859, n_860, n_861, n_862, n_863, n_864, n_865;
  wire n_866, n_867, n_868, n_869, n_870, n_871, n_872, n_873;
  wire n_874, n_875, n_876, n_877, n_878, n_879, n_880, n_881;
  wire n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889;
  wire n_890, n_891, n_892, n_893, n_894, n_895, n_896, n_897;
  wire n_898, n_899, n_900, n_901, n_902, n_903, n_904, n_905;
  wire n_906, n_907, n_908, n_909, n_910, n_911, n_912, n_913;
  wire n_914, n_915, n_916, n_917, n_918, n_919, n_920, n_921;
  wire n_922, n_923, n_924, n_925, n_926, n_927, n_928, n_929;
  wire n_930, n_931, n_932, n_933, n_934, n_935, n_936, n_937;
  wire n_938, n_939, n_940, n_941, n_942, n_943, n_944, n_945;
  wire n_946, n_947, n_948, n_949, n_950, n_951, n_952, n_953;
  wire n_954, n_955, n_956, n_957, n_958, n_959, n_960, n_961;
  wire n_962, n_963, n_964, n_965, n_966, n_967, n_968, n_969;
  wire n_970, n_971, n_972, n_973, n_974, n_975, n_976, n_977;
  wire n_978, n_979, n_980, n_981, n_982, n_983, n_984, n_985;
  wire n_986, n_987;
  xor g1 (n_831, A[0], B[0]);
  nand g2 (n_194, A[0], B[0]);
  nand g3 (n_195, A[0], CI);
  nand g4 (n_196, B[0], CI);
  nand g5 (n_198, n_194, n_195, n_196);
  nor g6 (n_197, A[1], B[1]);
  nand g7 (n_200, A[1], B[1]);
  nor g8 (n_207, A[2], B[2]);
  nand g9 (n_202, A[2], B[2]);
  nor g10 (n_203, A[3], B[3]);
  nand g11 (n_204, A[3], B[3]);
  nor g12 (n_213, A[4], B[4]);
  nand g13 (n_208, A[4], B[4]);
  nor g14 (n_209, A[5], B[5]);
  nand g15 (n_210, A[5], B[5]);
  nor g16 (n_219, A[6], B[6]);
  nand g17 (n_214, A[6], B[6]);
  nor g18 (n_215, A[7], B[7]);
  nand g19 (n_216, A[7], B[7]);
  nor g20 (n_225, A[8], B[8]);
  nand g21 (n_220, A[8], B[8]);
  nor g22 (n_221, A[9], B[9]);
  nand g23 (n_222, A[9], B[9]);
  nor g24 (n_231, A[10], B[10]);
  nand g25 (n_226, A[10], B[10]);
  nor g26 (n_227, A[11], B[11]);
  nand g27 (n_228, A[11], B[11]);
  nor g28 (n_237, A[12], B[12]);
  nand g29 (n_232, A[12], B[12]);
  nor g30 (n_233, A[13], B[13]);
  nand g31 (n_234, A[13], B[13]);
  nor g32 (n_243, A[14], B[14]);
  nand g33 (n_238, A[14], B[14]);
  nor g34 (n_239, A[15], B[15]);
  nand g35 (n_240, A[15], B[15]);
  nor g36 (n_249, A[16], B[16]);
  nand g37 (n_244, A[16], B[16]);
  nor g38 (n_245, A[17], B[17]);
  nand g39 (n_246, A[17], B[17]);
  nor g40 (n_255, A[18], B[18]);
  nand g41 (n_250, A[18], B[18]);
  nor g42 (n_251, A[19], B[19]);
  nand g43 (n_252, A[19], B[19]);
  nor g44 (n_261, A[20], B[20]);
  nand g45 (n_256, A[20], B[20]);
  nor g46 (n_257, A[21], B[21]);
  nand g47 (n_258, A[21], B[21]);
  nor g48 (n_267, A[22], B[22]);
  nand g49 (n_262, A[22], B[22]);
  nor g50 (n_263, A[23], B[23]);
  nand g51 (n_264, A[23], B[23]);
  nor g52 (n_273, A[24], B[24]);
  nand g53 (n_268, A[24], B[24]);
  nor g54 (n_269, A[25], B[25]);
  nand g55 (n_270, A[25], B[25]);
  nor g56 (n_279, A[26], B[26]);
  nand g57 (n_274, A[26], B[26]);
  nor g58 (n_275, A[27], B[27]);
  nand g59 (n_276, A[27], B[27]);
  nor g60 (n_285, A[28], B[28]);
  nand g61 (n_280, A[28], B[28]);
  nor g62 (n_281, A[29], B[29]);
  nand g63 (n_282, A[29], B[29]);
  nor g64 (n_291, A[30], B[30]);
  nand g65 (n_286, A[30], B[30]);
  nor g66 (n_287, A[31], B[31]);
  nand g67 (n_288, A[31], B[31]);
  nor g68 (n_297, A[32], B[32]);
  nand g69 (n_292, A[32], B[32]);
  nor g70 (n_293, A[33], B[33]);
  nand g71 (n_294, A[33], B[33]);
  nor g72 (n_303, A[34], B[34]);
  nand g73 (n_298, A[34], B[34]);
  nor g74 (n_299, A[35], B[35]);
  nand g75 (n_300, A[35], B[35]);
  nor g76 (n_309, A[36], B[36]);
  nand g77 (n_304, A[36], B[36]);
  nor g78 (n_305, A[37], B[37]);
  nand g79 (n_306, A[37], B[37]);
  nor g80 (n_315, A[38], B[38]);
  nand g81 (n_310, A[38], B[38]);
  nor g82 (n_311, A[39], B[39]);
  nand g83 (n_312, A[39], B[39]);
  nor g84 (n_321, A[40], B[40]);
  nand g85 (n_316, A[40], B[40]);
  nor g86 (n_317, A[41], B[41]);
  nand g87 (n_318, A[41], B[41]);
  nor g88 (n_327, A[42], B[42]);
  nand g89 (n_322, A[42], B[42]);
  nor g90 (n_323, A[43], B[43]);
  nand g91 (n_324, A[43], B[43]);
  nor g92 (n_333, A[44], B[44]);
  nand g93 (n_328, A[44], B[44]);
  nor g94 (n_329, A[45], B[45]);
  nand g95 (n_330, A[45], B[45]);
  nor g96 (n_339, A[46], B[46]);
  nand g97 (n_334, A[46], B[46]);
  nor g98 (n_335, A[47], B[47]);
  nand g99 (n_336, A[47], B[47]);
  nor g100 (n_345, A[48], B[48]);
  nand g101 (n_340, A[48], B[48]);
  nor g102 (n_341, A[49], B[49]);
  nand g103 (n_342, A[49], B[49]);
  nor g104 (n_351, A[50], B[50]);
  nand g105 (n_346, A[50], B[50]);
  nor g106 (n_347, A[51], B[51]);
  nand g107 (n_348, A[51], B[51]);
  nor g108 (n_357, A[52], B[52]);
  nand g109 (n_352, A[52], B[52]);
  nor g110 (n_353, A[53], B[53]);
  nand g111 (n_354, A[53], B[53]);
  nor g112 (n_363, A[54], B[54]);
  nand g113 (n_358, A[54], B[54]);
  nor g114 (n_359, A[55], B[55]);
  nand g115 (n_360, A[55], B[55]);
  nor g116 (n_369, A[56], B[56]);
  nand g117 (n_364, A[56], B[56]);
  nor g118 (n_365, A[57], B[57]);
  nand g119 (n_366, A[57], B[57]);
  nor g120 (n_375, A[58], B[58]);
  nand g121 (n_370, A[58], B[58]);
  nor g122 (n_371, A[59], B[59]);
  nand g123 (n_372, A[59], B[59]);
  nor g124 (n_381, A[60], B[60]);
  nand g125 (n_376, A[60], B[60]);
  nor g126 (n_377, A[61], B[61]);
  nand g127 (n_378, A[61], B[61]);
  nor g128 (n_387, A[62], B[62]);
  nand g129 (n_382, A[62], B[62]);
  nor g130 (n_383, A[63], B[63]);
  nand g131 (n_384, A[63], B[63]);
  nand g134 (n_389, n_200, n_837);
  nor g135 (n_205, n_202, n_203);
  nor g138 (n_388, n_207, n_203);
  nor g139 (n_211, n_208, n_209);
  nor g142 (n_398, n_213, n_209);
  nor g143 (n_217, n_214, n_215);
  nor g146 (n_392, n_219, n_215);
  nor g147 (n_223, n_220, n_221);
  nor g150 (n_405, n_225, n_221);
  nor g151 (n_229, n_226, n_227);
  nor g154 (n_399, n_231, n_227);
  nor g155 (n_235, n_232, n_233);
  nor g158 (n_412, n_237, n_233);
  nor g159 (n_241, n_238, n_239);
  nor g162 (n_406, n_243, n_239);
  nor g163 (n_247, n_244, n_245);
  nor g166 (n_419, n_249, n_245);
  nor g167 (n_253, n_250, n_251);
  nor g170 (n_413, n_255, n_251);
  nor g171 (n_259, n_256, n_257);
  nor g174 (n_426, n_261, n_257);
  nor g175 (n_265, n_262, n_263);
  nor g178 (n_420, n_267, n_263);
  nor g179 (n_271, n_268, n_269);
  nor g182 (n_433, n_273, n_269);
  nor g183 (n_277, n_274, n_275);
  nor g186 (n_427, n_279, n_275);
  nor g187 (n_283, n_280, n_281);
  nor g190 (n_440, n_285, n_281);
  nor g191 (n_289, n_286, n_287);
  nor g194 (n_434, n_291, n_287);
  nor g195 (n_295, n_292, n_293);
  nor g198 (n_447, n_297, n_293);
  nor g199 (n_301, n_298, n_299);
  nor g202 (n_441, n_303, n_299);
  nor g203 (n_307, n_304, n_305);
  nor g206 (n_454, n_309, n_305);
  nor g207 (n_313, n_310, n_311);
  nor g210 (n_448, n_315, n_311);
  nor g211 (n_319, n_316, n_317);
  nor g214 (n_461, n_321, n_317);
  nor g215 (n_325, n_322, n_323);
  nor g218 (n_455, n_327, n_323);
  nor g219 (n_331, n_328, n_329);
  nor g222 (n_468, n_333, n_329);
  nor g223 (n_337, n_334, n_335);
  nor g226 (n_462, n_339, n_335);
  nor g227 (n_343, n_340, n_341);
  nor g230 (n_475, n_345, n_341);
  nor g231 (n_349, n_346, n_347);
  nor g234 (n_469, n_351, n_347);
  nor g235 (n_355, n_352, n_353);
  nor g238 (n_482, n_357, n_353);
  nor g239 (n_361, n_358, n_359);
  nor g242 (n_476, n_363, n_359);
  nor g243 (n_367, n_364, n_365);
  nor g246 (n_489, n_369, n_365);
  nor g247 (n_373, n_370, n_371);
  nor g250 (n_483, n_375, n_371);
  nor g251 (n_379, n_376, n_377);
  nor g254 (n_496, n_381, n_377);
  nand g259 (n_391, n_388, n_389);
  nand g260 (n_498, n_838, n_391);
  nand g265 (n_497, n_398, n_392);
  nand g270 (n_507, n_405, n_399);
  nand g275 (n_502, n_412, n_406);
  nand g280 (n_513, n_419, n_413);
  nand g285 (n_508, n_426, n_420);
  nand g290 (n_519, n_433, n_427);
  nand g295 (n_514, n_440, n_434);
  nand g300 (n_525, n_447, n_441);
  nand g305 (n_520, n_454, n_448);
  nand g310 (n_531, n_461, n_455);
  nand g315 (n_526, n_468, n_462);
  nand g320 (n_537, n_475, n_469);
  nand g325 (n_532, n_482, n_476);
  nand g330 (n_543, n_489, n_483);
  nand g338 (n_545, n_931, n_940);
  nor g339 (n_505, n_502, n_503);
  nor g342 (n_544, n_507, n_502);
  nor g343 (n_511, n_508, n_509);
  nor g346 (n_554, n_513, n_508);
  nor g347 (n_517, n_514, n_515);
  nor g350 (n_548, n_519, n_514);
  nor g351 (n_523, n_520, n_521);
  nor g354 (n_561, n_525, n_520);
  nor g355 (n_529, n_526, n_527);
  nor g358 (n_555, n_531, n_526);
  nor g359 (n_535, n_532, n_533);
  nor g362 (n_568, n_537, n_532);
  nand g367 (n_547, n_544, n_545);
  nand g368 (n_570, n_941, n_547);
  nand g373 (n_569, n_554, n_548);
  nand g378 (n_579, n_561, n_555);
  nand g386 (n_581, n_948, n_953);
  nand g395 (n_588, n_949, n_958);
  nand g396 (n_586, n_554, n_570);
  nand g397 (n_594, n_549, n_586);
  nand g398 (n_587, n_561, n_581);
  nand g399 (n_599, n_556, n_587);
  nand g400 (n_589, n_568, n_588);
  nand g401 (n_604, n_944, n_589);
  nand g404 (n_609, n_503, n_950);
  nand g407 (n_612, n_509, n_954);
  nand g410 (n_615, n_515, n_959);
  nand g413 (n_618, n_521, n_960);
  nand g416 (n_621, n_527, n_966);
  nand g419 (n_624, n_533, n_967);
  nand g422 (n_627, n_938, n_975);
  nand g423 (n_607, n_398, n_498);
  nand g424 (n_633, n_393, n_607);
  nand g425 (n_608, n_405, n_545);
  nand g426 (n_638, n_400, n_608);
  nand g427 (n_610, n_412, n_609);
  nand g428 (n_643, n_407, n_610);
  nand g429 (n_611, n_419, n_570);
  nand g430 (n_648, n_414, n_611);
  nand g431 (n_613, n_426, n_612);
  nand g432 (n_653, n_421, n_613);
  nand g433 (n_614, n_433, n_594);
  nand g434 (n_658, n_428, n_614);
  nand g435 (n_616, n_440, n_615);
  nand g436 (n_663, n_435, n_616);
  nand g437 (n_617, n_447, n_581);
  nand g438 (n_668, n_442, n_617);
  nand g439 (n_619, n_454, n_618);
  nand g440 (n_673, n_449, n_619);
  nand g441 (n_620, n_461, n_599);
  nand g442 (n_678, n_456, n_620);
  nand g443 (n_622, n_468, n_621);
  nand g444 (n_683, n_463, n_622);
  nand g445 (n_623, n_475, n_588);
  nand g446 (n_688, n_470, n_623);
  nand g447 (n_625, n_482, n_624);
  nand g448 (n_693, n_477, n_625);
  nand g449 (n_626, n_489, n_604);
  nand g450 (n_698, n_484, n_626);
  nand g451 (n_628, n_496, n_627);
  nand g452 (n_703, n_853, n_628);
  nand g455 (n_709, n_202, n_939);
  nand g458 (n_713, n_208, n_945);
  nand g461 (n_717, n_214, n_951);
  nand g464 (n_721, n_220, n_952);
  nand g467 (n_725, n_226, n_955);
  nand g470 (n_729, n_232, n_956);
  nand g473 (n_733, n_238, n_961);
  nand g476 (n_737, n_244, n_957);
  nand g479 (n_741, n_250, n_962);
  nand g482 (n_745, n_256, n_963);
  nand g485 (n_749, n_262, n_968);
  nand g488 (n_753, n_268, n_964);
  nand g491 (n_757, n_274, n_969);
  nand g494 (n_761, n_280, n_970);
  nand g497 (n_765, n_286, n_976);
  nand g500 (n_769, n_292, n_965);
  nand g503 (n_773, n_298, n_971);
  nand g506 (n_777, n_304, n_972);
  nand g509 (n_781, n_310, n_977);
  nand g512 (n_785, n_316, n_973);
  nand g515 (n_789, n_322, n_978);
  nand g518 (n_793, n_328, n_979);
  nand g521 (n_797, n_334, n_983);
  nand g524 (n_801, n_340, n_974);
  nand g527 (n_805, n_346, n_980);
  nand g530 (n_809, n_352, n_981);
  nand g533 (n_813, n_358, n_984);
  nand g536 (n_817, n_364, n_982);
  nand g539 (n_821, n_370, n_985);
  nand g542 (n_825, n_376, n_986);
  nand g545 (n_829, n_382, n_987);
  xnor g547 (Z[1], n_198, n_854);
  xnor g549 (Z[2], n_389, n_855);
  xnor g552 (Z[3], n_709, n_856);
  xnor g554 (Z[4], n_498, n_857);
  xnor g557 (Z[5], n_713, n_858);
  xnor g559 (Z[6], n_633, n_859);
  xnor g562 (Z[7], n_717, n_860);
  xnor g564 (Z[8], n_545, n_861);
  xnor g567 (Z[9], n_721, n_862);
  xnor g569 (Z[10], n_638, n_863);
  xnor g572 (Z[11], n_725, n_864);
  xnor g574 (Z[12], n_609, n_865);
  xnor g577 (Z[13], n_729, n_866);
  xnor g579 (Z[14], n_643, n_867);
  xnor g582 (Z[15], n_733, n_868);
  xnor g584 (Z[16], n_570, n_869);
  xnor g587 (Z[17], n_737, n_870);
  xnor g589 (Z[18], n_648, n_871);
  xnor g592 (Z[19], n_741, n_872);
  xnor g594 (Z[20], n_612, n_873);
  xnor g597 (Z[21], n_745, n_874);
  xnor g599 (Z[22], n_653, n_875);
  xnor g602 (Z[23], n_749, n_876);
  xnor g604 (Z[24], n_594, n_877);
  xnor g607 (Z[25], n_753, n_878);
  xnor g609 (Z[26], n_658, n_879);
  xnor g612 (Z[27], n_757, n_880);
  xnor g614 (Z[28], n_615, n_881);
  xnor g617 (Z[29], n_761, n_882);
  xnor g619 (Z[30], n_663, n_883);
  xnor g622 (Z[31], n_765, n_884);
  xnor g624 (Z[32], n_581, n_885);
  xnor g627 (Z[33], n_769, n_886);
  xnor g629 (Z[34], n_668, n_887);
  xnor g632 (Z[35], n_773, n_888);
  xnor g634 (Z[36], n_618, n_889);
  xnor g637 (Z[37], n_777, n_890);
  xnor g639 (Z[38], n_673, n_891);
  xnor g642 (Z[39], n_781, n_892);
  xnor g644 (Z[40], n_599, n_893);
  xnor g647 (Z[41], n_785, n_894);
  xnor g649 (Z[42], n_678, n_895);
  xnor g652 (Z[43], n_789, n_896);
  xnor g654 (Z[44], n_621, n_897);
  xnor g657 (Z[45], n_793, n_898);
  xnor g659 (Z[46], n_683, n_899);
  xnor g662 (Z[47], n_797, n_900);
  xnor g664 (Z[48], n_588, n_901);
  xnor g667 (Z[49], n_801, n_902);
  xnor g669 (Z[50], n_688, n_903);
  xnor g672 (Z[51], n_805, n_904);
  xnor g674 (Z[52], n_624, n_905);
  xnor g677 (Z[53], n_809, n_906);
  xnor g679 (Z[54], n_693, n_907);
  xnor g682 (Z[55], n_813, n_908);
  xnor g684 (Z[56], n_604, n_909);
  xnor g687 (Z[57], n_817, n_910);
  xnor g689 (Z[58], n_698, n_911);
  xnor g692 (Z[59], n_821, n_912);
  xnor g694 (Z[60], n_627, n_913);
  xnor g697 (Z[61], n_825, n_914);
  xnor g699 (Z[62], n_703, n_915);
  xnor g702 (Z[63], n_829, n_916);
  xor g703 (Z[0], CI, n_831);
  or g704 (n_837, n_197, wc);
  not gc (wc, n_198);
  and g705 (n_838, wc0, n_204);
  not gc0 (wc0, n_205);
  and g706 (n_393, wc1, n_210);
  not gc1 (wc1, n_211);
  and g707 (n_839, wc2, n_216);
  not gc2 (wc2, n_217);
  and g708 (n_400, wc3, n_222);
  not gc3 (wc3, n_223);
  and g709 (n_840, wc4, n_228);
  not gc4 (wc4, n_229);
  and g710 (n_407, wc5, n_234);
  not gc5 (wc5, n_235);
  and g711 (n_841, wc6, n_240);
  not gc6 (wc6, n_241);
  and g712 (n_414, wc7, n_246);
  not gc7 (wc7, n_247);
  and g713 (n_842, wc8, n_252);
  not gc8 (wc8, n_253);
  and g714 (n_421, wc9, n_258);
  not gc9 (wc9, n_259);
  and g715 (n_843, wc10, n_264);
  not gc10 (wc10, n_265);
  and g716 (n_428, wc11, n_270);
  not gc11 (wc11, n_271);
  and g717 (n_844, wc12, n_276);
  not gc12 (wc12, n_277);
  and g718 (n_435, wc13, n_282);
  not gc13 (wc13, n_283);
  and g719 (n_845, wc14, n_288);
  not gc14 (wc14, n_289);
  and g720 (n_442, wc15, n_294);
  not gc15 (wc15, n_295);
  and g721 (n_846, wc16, n_300);
  not gc16 (wc16, n_301);
  and g722 (n_449, wc17, n_306);
  not gc17 (wc17, n_307);
  and g723 (n_847, wc18, n_312);
  not gc18 (wc18, n_313);
  and g724 (n_456, wc19, n_318);
  not gc19 (wc19, n_319);
  and g725 (n_848, wc20, n_324);
  not gc20 (wc20, n_325);
  and g726 (n_463, wc21, n_330);
  not gc21 (wc21, n_331);
  and g727 (n_849, wc22, n_336);
  not gc22 (wc22, n_337);
  and g728 (n_470, wc23, n_342);
  not gc23 (wc23, n_343);
  and g729 (n_850, wc24, n_348);
  not gc24 (wc24, n_349);
  and g730 (n_477, wc25, n_354);
  not gc25 (wc25, n_355);
  and g731 (n_851, wc26, n_360);
  not gc26 (wc26, n_361);
  and g732 (n_484, wc27, n_366);
  not gc27 (wc27, n_367);
  and g733 (n_852, wc28, n_372);
  not gc28 (wc28, n_373);
  and g734 (n_853, wc29, n_378);
  not gc29 (wc29, n_379);
  or g735 (n_854, wc30, n_197);
  not gc30 (wc30, n_200);
  or g736 (n_855, wc31, n_207);
  not gc31 (wc31, n_202);
  or g737 (n_856, wc32, n_203);
  not gc32 (wc32, n_204);
  or g738 (n_857, wc33, n_213);
  not gc33 (wc33, n_208);
  or g739 (n_858, wc34, n_209);
  not gc34 (wc34, n_210);
  or g740 (n_859, wc35, n_219);
  not gc35 (wc35, n_214);
  or g741 (n_860, wc36, n_215);
  not gc36 (wc36, n_216);
  or g742 (n_861, wc37, n_225);
  not gc37 (wc37, n_220);
  or g743 (n_862, wc38, n_221);
  not gc38 (wc38, n_222);
  or g744 (n_863, wc39, n_231);
  not gc39 (wc39, n_226);
  or g745 (n_864, wc40, n_227);
  not gc40 (wc40, n_228);
  or g746 (n_865, wc41, n_237);
  not gc41 (wc41, n_232);
  or g747 (n_866, wc42, n_233);
  not gc42 (wc42, n_234);
  or g748 (n_867, wc43, n_243);
  not gc43 (wc43, n_238);
  or g749 (n_868, wc44, n_239);
  not gc44 (wc44, n_240);
  or g750 (n_869, wc45, n_249);
  not gc45 (wc45, n_244);
  or g751 (n_870, wc46, n_245);
  not gc46 (wc46, n_246);
  or g752 (n_871, wc47, n_255);
  not gc47 (wc47, n_250);
  or g753 (n_872, wc48, n_251);
  not gc48 (wc48, n_252);
  or g754 (n_873, wc49, n_261);
  not gc49 (wc49, n_256);
  or g755 (n_874, wc50, n_257);
  not gc50 (wc50, n_258);
  or g756 (n_875, wc51, n_267);
  not gc51 (wc51, n_262);
  or g757 (n_876, wc52, n_263);
  not gc52 (wc52, n_264);
  or g758 (n_877, wc53, n_273);
  not gc53 (wc53, n_268);
  or g759 (n_878, wc54, n_269);
  not gc54 (wc54, n_270);
  or g760 (n_879, wc55, n_279);
  not gc55 (wc55, n_274);
  or g761 (n_880, wc56, n_275);
  not gc56 (wc56, n_276);
  or g762 (n_881, wc57, n_285);
  not gc57 (wc57, n_280);
  or g763 (n_882, wc58, n_281);
  not gc58 (wc58, n_282);
  or g764 (n_883, wc59, n_291);
  not gc59 (wc59, n_286);
  or g765 (n_884, wc60, n_287);
  not gc60 (wc60, n_288);
  or g766 (n_885, wc61, n_297);
  not gc61 (wc61, n_292);
  or g767 (n_886, wc62, n_293);
  not gc62 (wc62, n_294);
  or g768 (n_887, wc63, n_303);
  not gc63 (wc63, n_298);
  or g769 (n_888, wc64, n_299);
  not gc64 (wc64, n_300);
  or g770 (n_889, wc65, n_309);
  not gc65 (wc65, n_304);
  or g771 (n_890, wc66, n_305);
  not gc66 (wc66, n_306);
  or g772 (n_891, wc67, n_315);
  not gc67 (wc67, n_310);
  or g773 (n_892, wc68, n_311);
  not gc68 (wc68, n_312);
  or g774 (n_893, wc69, n_321);
  not gc69 (wc69, n_316);
  or g775 (n_894, wc70, n_317);
  not gc70 (wc70, n_318);
  or g776 (n_895, wc71, n_327);
  not gc71 (wc71, n_322);
  or g777 (n_896, wc72, n_323);
  not gc72 (wc72, n_324);
  or g778 (n_897, wc73, n_333);
  not gc73 (wc73, n_328);
  or g779 (n_898, wc74, n_329);
  not gc74 (wc74, n_330);
  or g780 (n_899, wc75, n_339);
  not gc75 (wc75, n_334);
  or g781 (n_900, wc76, n_335);
  not gc76 (wc76, n_336);
  or g782 (n_901, wc77, n_345);
  not gc77 (wc77, n_340);
  or g783 (n_902, wc78, n_341);
  not gc78 (wc78, n_342);
  or g784 (n_903, wc79, n_351);
  not gc79 (wc79, n_346);
  or g785 (n_904, wc80, n_347);
  not gc80 (wc80, n_348);
  or g786 (n_905, wc81, n_357);
  not gc81 (wc81, n_352);
  or g787 (n_906, wc82, n_353);
  not gc82 (wc82, n_354);
  or g788 (n_907, wc83, n_363);
  not gc83 (wc83, n_358);
  or g789 (n_908, wc84, n_359);
  not gc84 (wc84, n_360);
  or g790 (n_909, wc85, n_369);
  not gc85 (wc85, n_364);
  or g791 (n_910, wc86, n_365);
  not gc86 (wc86, n_366);
  or g792 (n_911, wc87, n_375);
  not gc87 (wc87, n_370);
  or g793 (n_912, wc88, n_371);
  not gc88 (wc88, n_372);
  or g794 (n_913, wc89, n_381);
  not gc89 (wc89, n_376);
  or g795 (n_914, wc90, n_377);
  not gc90 (wc90, n_378);
  or g796 (n_915, wc91, n_387);
  not gc91 (wc91, n_382);
  or g797 (n_916, wc92, n_383);
  not gc92 (wc92, n_384);
  and g798 (n_917, wc93, n_392);
  not gc93 (wc93, n_393);
  and g799 (n_918, wc94, n_399);
  not gc94 (wc94, n_400);
  and g800 (n_919, wc95, n_406);
  not gc95 (wc95, n_407);
  and g801 (n_920, wc96, n_413);
  not gc96 (wc96, n_414);
  and g802 (n_921, wc97, n_420);
  not gc97 (wc97, n_421);
  and g803 (n_922, wc98, n_427);
  not gc98 (wc98, n_428);
  and g804 (n_923, wc99, n_434);
  not gc99 (wc99, n_435);
  and g805 (n_924, wc100, n_441);
  not gc100 (wc100, n_442);
  and g806 (n_925, wc101, n_448);
  not gc101 (wc101, n_449);
  and g807 (n_926, wc102, n_455);
  not gc102 (wc102, n_456);
  and g808 (n_927, wc103, n_462);
  not gc103 (wc103, n_463);
  and g809 (n_928, wc104, n_469);
  not gc104 (wc104, n_470);
  and g810 (n_929, wc105, n_476);
  not gc105 (wc105, n_477);
  and g811 (n_930, wc106, n_483);
  not gc106 (wc106, n_484);
  and g812 (n_931, wc107, n_839);
  not gc107 (wc107, n_917);
  and g813 (n_503, wc108, n_840);
  not gc108 (wc108, n_918);
  and g814 (n_932, wc109, n_841);
  not gc109 (wc109, n_919);
  and g815 (n_509, wc110, n_842);
  not gc110 (wc110, n_920);
  and g816 (n_933, wc111, n_843);
  not gc111 (wc111, n_921);
  and g817 (n_515, wc112, n_844);
  not gc112 (wc112, n_922);
  and g818 (n_934, wc113, n_845);
  not gc113 (wc113, n_923);
  and g819 (n_521, wc114, n_846);
  not gc114 (wc114, n_924);
  and g820 (n_935, wc115, n_847);
  not gc115 (wc115, n_925);
  and g821 (n_527, wc116, n_848);
  not gc116 (wc116, n_926);
  and g822 (n_936, wc117, n_849);
  not gc117 (wc117, n_927);
  and g823 (n_533, wc118, n_850);
  not gc118 (wc118, n_928);
  and g824 (n_937, wc119, n_851);
  not gc119 (wc119, n_929);
  and g825 (n_938, wc120, n_852);
  not gc120 (wc120, n_930);
  or g826 (n_939, wc121, n_207);
  not gc121 (wc121, n_389);
  or g827 (n_940, n_497, wc122);
  not gc122 (wc122, n_498);
  and g828 (n_941, n_932, wc123);
  not gc123 (wc123, n_505);
  and g829 (n_549, n_933, wc124);
  not gc124 (wc124, n_511);
  and g830 (n_942, n_934, wc125);
  not gc125 (wc125, n_517);
  and g831 (n_556, n_935, wc126);
  not gc126 (wc126, n_523);
  and g832 (n_943, n_936, wc127);
  not gc127 (wc127, n_529);
  and g833 (n_944, n_937, wc128);
  not gc128 (wc128, n_535);
  or g834 (n_945, wc129, n_213);
  not gc129 (wc129, n_498);
  and g835 (n_946, wc130, n_548);
  not gc130 (wc130, n_549);
  and g836 (n_947, wc131, n_555);
  not gc131 (wc131, n_556);
  and g837 (n_948, wc132, n_942);
  not gc132 (wc132, n_946);
  and g838 (n_949, wc133, n_943);
  not gc133 (wc133, n_947);
  or g839 (n_950, wc134, n_507);
  not gc134 (wc134, n_545);
  or g840 (n_951, wc135, n_219);
  not gc135 (wc135, n_633);
  or g841 (n_952, wc136, n_225);
  not gc136 (wc136, n_545);
  or g842 (n_953, n_569, wc137);
  not gc137 (wc137, n_570);
  or g843 (n_954, wc138, n_513);
  not gc138 (wc138, n_570);
  or g844 (n_955, wc139, n_231);
  not gc139 (wc139, n_638);
  or g845 (n_956, wc140, n_237);
  not gc140 (wc140, n_609);
  or g846 (n_957, wc141, n_249);
  not gc141 (wc141, n_570);
  or g847 (n_958, wc142, n_579);
  not gc142 (wc142, n_581);
  or g848 (n_959, wc143, n_519);
  not gc143 (wc143, n_594);
  or g849 (n_960, wc144, n_525);
  not gc144 (wc144, n_581);
  or g850 (n_961, wc145, n_243);
  not gc145 (wc145, n_643);
  or g851 (n_962, wc146, n_255);
  not gc146 (wc146, n_648);
  or g852 (n_963, wc147, n_261);
  not gc147 (wc147, n_612);
  or g853 (n_964, wc148, n_273);
  not gc148 (wc148, n_594);
  or g854 (n_965, wc149, n_297);
  not gc149 (wc149, n_581);
  or g855 (n_966, wc150, n_531);
  not gc150 (wc150, n_599);
  or g856 (n_967, wc151, n_537);
  not gc151 (wc151, n_588);
  or g857 (n_968, wc152, n_267);
  not gc152 (wc152, n_653);
  or g858 (n_969, wc153, n_279);
  not gc153 (wc153, n_658);
  or g859 (n_970, wc154, n_285);
  not gc154 (wc154, n_615);
  or g860 (n_971, wc155, n_303);
  not gc155 (wc155, n_668);
  or g861 (n_972, wc156, n_309);
  not gc156 (wc156, n_618);
  or g862 (n_973, wc157, n_321);
  not gc157 (wc157, n_599);
  or g863 (n_974, wc158, n_345);
  not gc158 (wc158, n_588);
  or g864 (n_975, wc159, n_543);
  not gc159 (wc159, n_604);
  or g865 (n_976, wc160, n_291);
  not gc160 (wc160, n_663);
  or g866 (n_977, wc161, n_315);
  not gc161 (wc161, n_673);
  or g867 (n_978, wc162, n_327);
  not gc162 (wc162, n_678);
  or g868 (n_979, wc163, n_333);
  not gc163 (wc163, n_621);
  or g869 (n_980, wc164, n_351);
  not gc164 (wc164, n_688);
  or g870 (n_981, wc165, n_357);
  not gc165 (wc165, n_624);
  or g871 (n_982, wc166, n_369);
  not gc166 (wc166, n_604);
  or g872 (n_983, wc167, n_339);
  not gc167 (wc167, n_683);
  or g873 (n_984, wc168, n_363);
  not gc168 (wc168, n_693);
  or g874 (n_985, wc169, n_375);
  not gc169 (wc169, n_698);
  or g875 (n_986, wc170, n_381);
  not gc170 (wc170, n_627);
  or g876 (n_987, wc171, n_387);
  not gc171 (wc171, n_703);
endmodule

module add_unsigned_carry_2513_GENERIC(A, B, CI, Z);
  input [63:0] A, B;
  input CI;
  output [63:0] Z;
  wire [63:0] A, B;
  wire CI;
  wire [63:0] Z;
  add_unsigned_carry_2513_GENERIC_REAL g1(.A (A), .B (B), .CI (CI), .Z
       (Z));
endmodule

module add_unsigned_carry_2513_1_GENERIC_REAL(A, B, CI, Z);
// synthesis_equation add_unsigned_carry
  input [63:0] A, B;
  input CI;
  output [63:0] Z;
  wire [63:0] A, B;
  wire CI;
  wire [63:0] Z;
  wire n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201;
  wire n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209;
  wire n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225;
  wire n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241;
  wire n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249;
  wire n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257;
  wire n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265;
  wire n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273;
  wire n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281;
  wire n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289;
  wire n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297;
  wire n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313;
  wire n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329;
  wire n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345;
  wire n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353;
  wire n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361;
  wire n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369;
  wire n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377;
  wire n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385;
  wire n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393;
  wire n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401;
  wire n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409;
  wire n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417;
  wire n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425;
  wire n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433;
  wire n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457;
  wire n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465;
  wire n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473;
  wire n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481;
  wire n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489;
  wire n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497;
  wire n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505;
  wire n_506, n_507, n_508, n_512;
  nand g1 (n_194, A[0], B[0]);
  nand g2 (n_195, A[0], CI);
  nand g3 (n_196, B[0], CI);
  nand g4 (n_198, n_194, n_195, n_196);
  xor g5 (n_197, A[0], B[0]);
  xor g6 (Z[0], CI, n_197);
  nand g7 (n_199, A[1], B[1]);
  nand g8 (n_200, A[1], n_198);
  nand g9 (n_201, B[1], n_198);
  nand g10 (n_203, n_199, n_200, n_201);
  xor g11 (n_202, A[1], B[1]);
  xor g12 (Z[1], n_198, n_202);
  nand g13 (n_204, A[2], B[2]);
  nand g14 (n_205, A[2], n_203);
  nand g15 (n_206, B[2], n_203);
  nand g16 (n_208, n_204, n_205, n_206);
  xor g17 (n_207, A[2], B[2]);
  xor g18 (Z[2], n_203, n_207);
  nand g19 (n_209, A[3], B[3]);
  nand g20 (n_210, A[3], n_208);
  nand g21 (n_211, B[3], n_208);
  nand g22 (n_213, n_209, n_210, n_211);
  xor g23 (n_212, A[3], B[3]);
  xor g24 (Z[3], n_208, n_212);
  nand g25 (n_214, A[4], B[4]);
  nand g26 (n_215, A[4], n_213);
  nand g27 (n_216, B[4], n_213);
  nand g28 (n_218, n_214, n_215, n_216);
  xor g29 (n_217, A[4], B[4]);
  xor g30 (Z[4], n_213, n_217);
  nand g31 (n_219, A[5], B[5]);
  nand g32 (n_220, A[5], n_218);
  nand g33 (n_221, B[5], n_218);
  nand g34 (n_223, n_219, n_220, n_221);
  xor g35 (n_222, A[5], B[5]);
  xor g36 (Z[5], n_218, n_222);
  nand g37 (n_224, A[6], B[6]);
  nand g38 (n_225, A[6], n_223);
  nand g39 (n_226, B[6], n_223);
  nand g40 (n_228, n_224, n_225, n_226);
  xor g41 (n_227, A[6], B[6]);
  xor g42 (Z[6], n_223, n_227);
  nand g43 (n_229, A[7], B[7]);
  nand g44 (n_230, A[7], n_228);
  nand g45 (n_231, B[7], n_228);
  nand g46 (n_233, n_229, n_230, n_231);
  xor g47 (n_232, A[7], B[7]);
  xor g48 (Z[7], n_228, n_232);
  nand g49 (n_234, A[8], B[8]);
  nand g50 (n_235, A[8], n_233);
  nand g51 (n_236, B[8], n_233);
  nand g52 (n_238, n_234, n_235, n_236);
  xor g53 (n_237, A[8], B[8]);
  xor g54 (Z[8], n_233, n_237);
  nand g55 (n_239, A[9], B[9]);
  nand g56 (n_240, A[9], n_238);
  nand g57 (n_241, B[9], n_238);
  nand g58 (n_243, n_239, n_240, n_241);
  xor g59 (n_242, A[9], B[9]);
  xor g60 (Z[9], n_238, n_242);
  nand g61 (n_244, A[10], B[10]);
  nand g62 (n_245, A[10], n_243);
  nand g63 (n_246, B[10], n_243);
  nand g64 (n_248, n_244, n_245, n_246);
  xor g65 (n_247, A[10], B[10]);
  xor g66 (Z[10], n_243, n_247);
  nand g67 (n_249, A[11], B[11]);
  nand g68 (n_250, A[11], n_248);
  nand g69 (n_251, B[11], n_248);
  nand g70 (n_253, n_249, n_250, n_251);
  xor g71 (n_252, A[11], B[11]);
  xor g72 (Z[11], n_248, n_252);
  nand g73 (n_254, A[12], B[12]);
  nand g74 (n_255, A[12], n_253);
  nand g75 (n_256, B[12], n_253);
  nand g76 (n_258, n_254, n_255, n_256);
  xor g77 (n_257, A[12], B[12]);
  xor g78 (Z[12], n_253, n_257);
  nand g79 (n_259, A[13], B[13]);
  nand g80 (n_260, A[13], n_258);
  nand g81 (n_261, B[13], n_258);
  nand g82 (n_263, n_259, n_260, n_261);
  xor g83 (n_262, A[13], B[13]);
  xor g84 (Z[13], n_258, n_262);
  nand g85 (n_264, A[14], B[14]);
  nand g86 (n_265, A[14], n_263);
  nand g87 (n_266, B[14], n_263);
  nand g88 (n_268, n_264, n_265, n_266);
  xor g89 (n_267, A[14], B[14]);
  xor g90 (Z[14], n_263, n_267);
  nand g91 (n_269, A[15], B[15]);
  nand g92 (n_270, A[15], n_268);
  nand g93 (n_271, B[15], n_268);
  nand g94 (n_273, n_269, n_270, n_271);
  xor g95 (n_272, A[15], B[15]);
  xor g96 (Z[15], n_268, n_272);
  nand g97 (n_274, A[16], B[16]);
  nand g98 (n_275, A[16], n_273);
  nand g99 (n_276, B[16], n_273);
  nand g100 (n_278, n_274, n_275, n_276);
  xor g101 (n_277, A[16], B[16]);
  xor g102 (Z[16], n_273, n_277);
  nand g103 (n_279, A[17], B[17]);
  nand g104 (n_280, A[17], n_278);
  nand g105 (n_281, B[17], n_278);
  nand g106 (n_283, n_279, n_280, n_281);
  xor g107 (n_282, A[17], B[17]);
  xor g108 (Z[17], n_278, n_282);
  nand g109 (n_284, A[18], B[18]);
  nand g110 (n_285, A[18], n_283);
  nand g111 (n_286, B[18], n_283);
  nand g112 (n_288, n_284, n_285, n_286);
  xor g113 (n_287, A[18], B[18]);
  xor g114 (Z[18], n_283, n_287);
  nand g115 (n_289, A[19], B[19]);
  nand g116 (n_290, A[19], n_288);
  nand g117 (n_291, B[19], n_288);
  nand g118 (n_293, n_289, n_290, n_291);
  xor g119 (n_292, A[19], B[19]);
  xor g120 (Z[19], n_288, n_292);
  nand g121 (n_294, A[20], B[20]);
  nand g122 (n_295, A[20], n_293);
  nand g123 (n_296, B[20], n_293);
  nand g124 (n_298, n_294, n_295, n_296);
  xor g125 (n_297, A[20], B[20]);
  xor g126 (Z[20], n_293, n_297);
  nand g127 (n_299, A[21], B[21]);
  nand g128 (n_300, A[21], n_298);
  nand g129 (n_301, B[21], n_298);
  nand g130 (n_303, n_299, n_300, n_301);
  xor g131 (n_302, A[21], B[21]);
  xor g132 (Z[21], n_298, n_302);
  nand g133 (n_304, A[22], B[22]);
  nand g134 (n_305, A[22], n_303);
  nand g135 (n_306, B[22], n_303);
  nand g136 (n_308, n_304, n_305, n_306);
  xor g137 (n_307, A[22], B[22]);
  xor g138 (Z[22], n_303, n_307);
  nand g139 (n_309, A[23], B[23]);
  nand g140 (n_310, A[23], n_308);
  nand g141 (n_311, B[23], n_308);
  nand g142 (n_313, n_309, n_310, n_311);
  xor g143 (n_312, A[23], B[23]);
  xor g144 (Z[23], n_308, n_312);
  nand g145 (n_314, A[24], B[24]);
  nand g146 (n_315, A[24], n_313);
  nand g147 (n_316, B[24], n_313);
  nand g148 (n_318, n_314, n_315, n_316);
  xor g149 (n_317, A[24], B[24]);
  xor g150 (Z[24], n_313, n_317);
  nand g151 (n_319, A[25], B[25]);
  nand g152 (n_320, A[25], n_318);
  nand g153 (n_321, B[25], n_318);
  nand g154 (n_323, n_319, n_320, n_321);
  xor g155 (n_322, A[25], B[25]);
  xor g156 (Z[25], n_318, n_322);
  nand g157 (n_324, A[26], B[26]);
  nand g158 (n_325, A[26], n_323);
  nand g159 (n_326, B[26], n_323);
  nand g160 (n_328, n_324, n_325, n_326);
  xor g161 (n_327, A[26], B[26]);
  xor g162 (Z[26], n_323, n_327);
  nand g163 (n_329, A[27], B[27]);
  nand g164 (n_330, A[27], n_328);
  nand g165 (n_331, B[27], n_328);
  nand g166 (n_333, n_329, n_330, n_331);
  xor g167 (n_332, A[27], B[27]);
  xor g168 (Z[27], n_328, n_332);
  nand g169 (n_334, A[28], B[28]);
  nand g170 (n_335, A[28], n_333);
  nand g171 (n_336, B[28], n_333);
  nand g172 (n_338, n_334, n_335, n_336);
  xor g173 (n_337, A[28], B[28]);
  xor g174 (Z[28], n_333, n_337);
  nand g175 (n_339, A[29], B[29]);
  nand g176 (n_340, A[29], n_338);
  nand g177 (n_341, B[29], n_338);
  nand g178 (n_343, n_339, n_340, n_341);
  xor g179 (n_342, A[29], B[29]);
  xor g180 (Z[29], n_338, n_342);
  nand g181 (n_344, A[30], B[30]);
  nand g182 (n_345, A[30], n_343);
  nand g183 (n_346, B[30], n_343);
  nand g184 (n_348, n_344, n_345, n_346);
  xor g185 (n_347, A[30], B[30]);
  xor g186 (Z[30], n_343, n_347);
  nand g187 (n_349, A[31], B[31]);
  nand g188 (n_350, A[31], n_348);
  nand g189 (n_351, B[31], n_348);
  nand g190 (n_353, n_349, n_350, n_351);
  xor g191 (n_352, A[31], B[31]);
  xor g192 (Z[31], n_348, n_352);
  nand g193 (n_354, A[32], B[32]);
  nand g194 (n_355, A[32], n_353);
  nand g195 (n_356, B[32], n_353);
  nand g196 (n_358, n_354, n_355, n_356);
  xor g197 (n_357, A[32], B[32]);
  xor g198 (Z[32], n_353, n_357);
  nand g199 (n_359, A[33], B[33]);
  nand g200 (n_360, A[33], n_358);
  nand g201 (n_361, B[33], n_358);
  nand g202 (n_363, n_359, n_360, n_361);
  xor g203 (n_362, A[33], B[33]);
  xor g204 (Z[33], n_358, n_362);
  nand g205 (n_364, A[34], B[34]);
  nand g206 (n_365, A[34], n_363);
  nand g207 (n_366, B[34], n_363);
  nand g208 (n_368, n_364, n_365, n_366);
  xor g209 (n_367, A[34], B[34]);
  xor g210 (Z[34], n_363, n_367);
  nand g211 (n_369, A[35], B[35]);
  nand g212 (n_370, A[35], n_368);
  nand g213 (n_371, B[35], n_368);
  nand g214 (n_373, n_369, n_370, n_371);
  xor g215 (n_372, A[35], B[35]);
  xor g216 (Z[35], n_368, n_372);
  nand g217 (n_374, A[36], B[36]);
  nand g218 (n_375, A[36], n_373);
  nand g219 (n_376, B[36], n_373);
  nand g220 (n_378, n_374, n_375, n_376);
  xor g221 (n_377, A[36], B[36]);
  xor g222 (Z[36], n_373, n_377);
  nand g223 (n_379, A[37], B[37]);
  nand g224 (n_380, A[37], n_378);
  nand g225 (n_381, B[37], n_378);
  nand g226 (n_383, n_379, n_380, n_381);
  xor g227 (n_382, A[37], B[37]);
  xor g228 (Z[37], n_378, n_382);
  nand g229 (n_384, A[38], B[38]);
  nand g230 (n_385, A[38], n_383);
  nand g231 (n_386, B[38], n_383);
  nand g232 (n_388, n_384, n_385, n_386);
  xor g233 (n_387, A[38], B[38]);
  xor g234 (Z[38], n_383, n_387);
  nand g235 (n_389, A[39], B[39]);
  nand g236 (n_390, A[39], n_388);
  nand g237 (n_391, B[39], n_388);
  nand g238 (n_393, n_389, n_390, n_391);
  xor g239 (n_392, A[39], B[39]);
  xor g240 (Z[39], n_388, n_392);
  nand g241 (n_394, A[40], B[40]);
  nand g242 (n_395, A[40], n_393);
  nand g243 (n_396, B[40], n_393);
  nand g244 (n_398, n_394, n_395, n_396);
  xor g245 (n_397, A[40], B[40]);
  xor g246 (Z[40], n_393, n_397);
  nand g247 (n_399, A[41], B[41]);
  nand g248 (n_400, A[41], n_398);
  nand g249 (n_401, B[41], n_398);
  nand g250 (n_403, n_399, n_400, n_401);
  xor g251 (n_402, A[41], B[41]);
  xor g252 (Z[41], n_398, n_402);
  nand g253 (n_404, A[42], B[42]);
  nand g254 (n_405, A[42], n_403);
  nand g255 (n_406, B[42], n_403);
  nand g256 (n_408, n_404, n_405, n_406);
  xor g257 (n_407, A[42], B[42]);
  xor g258 (Z[42], n_403, n_407);
  nand g259 (n_409, A[43], B[43]);
  nand g260 (n_410, A[43], n_408);
  nand g261 (n_411, B[43], n_408);
  nand g262 (n_413, n_409, n_410, n_411);
  xor g263 (n_412, A[43], B[43]);
  xor g264 (Z[43], n_408, n_412);
  nand g265 (n_414, A[44], B[44]);
  nand g266 (n_415, A[44], n_413);
  nand g267 (n_416, B[44], n_413);
  nand g268 (n_418, n_414, n_415, n_416);
  xor g269 (n_417, A[44], B[44]);
  xor g270 (Z[44], n_413, n_417);
  nand g271 (n_419, A[45], B[45]);
  nand g272 (n_420, A[45], n_418);
  nand g273 (n_421, B[45], n_418);
  nand g274 (n_423, n_419, n_420, n_421);
  xor g275 (n_422, A[45], B[45]);
  xor g276 (Z[45], n_418, n_422);
  nand g277 (n_424, A[46], B[46]);
  nand g278 (n_425, A[46], n_423);
  nand g279 (n_426, B[46], n_423);
  nand g280 (n_428, n_424, n_425, n_426);
  xor g281 (n_427, A[46], B[46]);
  xor g282 (Z[46], n_423, n_427);
  nand g283 (n_429, A[47], B[47]);
  nand g284 (n_430, A[47], n_428);
  nand g285 (n_431, B[47], n_428);
  nand g286 (n_433, n_429, n_430, n_431);
  xor g287 (n_432, A[47], B[47]);
  xor g288 (Z[47], n_428, n_432);
  nand g289 (n_434, A[48], B[48]);
  nand g290 (n_435, A[48], n_433);
  nand g291 (n_436, B[48], n_433);
  nand g292 (n_438, n_434, n_435, n_436);
  xor g293 (n_437, A[48], B[48]);
  xor g294 (Z[48], n_433, n_437);
  nand g295 (n_439, A[49], B[49]);
  nand g296 (n_440, A[49], n_438);
  nand g297 (n_441, B[49], n_438);
  nand g298 (n_443, n_439, n_440, n_441);
  xor g299 (n_442, A[49], B[49]);
  xor g300 (Z[49], n_438, n_442);
  nand g301 (n_444, A[50], B[50]);
  nand g302 (n_445, A[50], n_443);
  nand g303 (n_446, B[50], n_443);
  nand g304 (n_448, n_444, n_445, n_446);
  xor g305 (n_447, A[50], B[50]);
  xor g306 (Z[50], n_443, n_447);
  nand g307 (n_449, A[51], B[51]);
  nand g308 (n_450, A[51], n_448);
  nand g309 (n_451, B[51], n_448);
  nand g310 (n_453, n_449, n_450, n_451);
  xor g311 (n_452, A[51], B[51]);
  xor g312 (Z[51], n_448, n_452);
  nand g313 (n_454, A[52], B[52]);
  nand g314 (n_455, A[52], n_453);
  nand g315 (n_456, B[52], n_453);
  nand g316 (n_458, n_454, n_455, n_456);
  xor g317 (n_457, A[52], B[52]);
  xor g318 (Z[52], n_453, n_457);
  nand g319 (n_459, A[53], B[53]);
  nand g320 (n_460, A[53], n_458);
  nand g321 (n_461, B[53], n_458);
  nand g322 (n_463, n_459, n_460, n_461);
  xor g323 (n_462, A[53], B[53]);
  xor g324 (Z[53], n_458, n_462);
  nand g325 (n_464, A[54], B[54]);
  nand g326 (n_465, A[54], n_463);
  nand g327 (n_466, B[54], n_463);
  nand g328 (n_468, n_464, n_465, n_466);
  xor g329 (n_467, A[54], B[54]);
  xor g330 (Z[54], n_463, n_467);
  nand g331 (n_469, A[55], B[55]);
  nand g332 (n_470, A[55], n_468);
  nand g333 (n_471, B[55], n_468);
  nand g334 (n_473, n_469, n_470, n_471);
  xor g335 (n_472, A[55], B[55]);
  xor g336 (Z[55], n_468, n_472);
  nand g337 (n_474, A[56], B[56]);
  nand g338 (n_475, A[56], n_473);
  nand g339 (n_476, B[56], n_473);
  nand g340 (n_478, n_474, n_475, n_476);
  xor g341 (n_477, A[56], B[56]);
  xor g342 (Z[56], n_473, n_477);
  nand g343 (n_479, A[57], B[57]);
  nand g344 (n_480, A[57], n_478);
  nand g345 (n_481, B[57], n_478);
  nand g346 (n_483, n_479, n_480, n_481);
  xor g347 (n_482, A[57], B[57]);
  xor g348 (Z[57], n_478, n_482);
  nand g349 (n_484, A[58], B[58]);
  nand g350 (n_485, A[58], n_483);
  nand g351 (n_486, B[58], n_483);
  nand g352 (n_488, n_484, n_485, n_486);
  xor g353 (n_487, A[58], B[58]);
  xor g354 (Z[58], n_483, n_487);
  nand g355 (n_489, A[59], B[59]);
  nand g356 (n_490, A[59], n_488);
  nand g357 (n_491, B[59], n_488);
  nand g358 (n_493, n_489, n_490, n_491);
  xor g359 (n_492, A[59], B[59]);
  xor g360 (Z[59], n_488, n_492);
  nand g361 (n_494, A[60], B[60]);
  nand g362 (n_495, A[60], n_493);
  nand g363 (n_496, B[60], n_493);
  nand g364 (n_498, n_494, n_495, n_496);
  xor g365 (n_497, A[60], B[60]);
  xor g366 (Z[60], n_493, n_497);
  nand g367 (n_499, A[61], B[61]);
  nand g368 (n_500, A[61], n_498);
  nand g369 (n_501, B[61], n_498);
  nand g370 (n_503, n_499, n_500, n_501);
  xor g371 (n_502, A[61], B[61]);
  xor g372 (Z[61], n_498, n_502);
  nand g373 (n_504, A[62], B[62]);
  nand g374 (n_505, A[62], n_503);
  nand g375 (n_506, B[62], n_503);
  nand g376 (n_508, n_504, n_505, n_506);
  xor g377 (n_507, A[62], B[62]);
  xor g378 (Z[62], n_503, n_507);
  xor g383 (n_512, A[63], B[63]);
  xor g384 (Z[63], n_508, n_512);
endmodule

module add_unsigned_carry_2513_1_GENERIC(A, B, CI, Z);
  input [63:0] A, B;
  input CI;
  output [63:0] Z;
  wire [63:0] A, B;
  wire CI;
  wire [63:0] Z;
  add_unsigned_carry_2513_1_GENERIC_REAL g1(.A (A), .B (B), .CI (CI),
       .Z (Z));
endmodule

module add_unsigned_carry_2520_GENERIC_REAL(A, B, CI, Z);
// synthesis_equation add_unsigned_carry
  input [54:0] A, B;
  input CI;
  output [54:0] Z;
  wire [54:0] A, B;
  wire CI;
  wire [54:0] Z;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190;
  wire n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198;
  wire n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206;
  wire n_207, n_208, n_209, n_210, n_211, n_212, n_213, n_214;
  wire n_215, n_216, n_217, n_218, n_219, n_220, n_221, n_222;
  wire n_223, n_224, n_225, n_226, n_227, n_228, n_229, n_230;
  wire n_231, n_232, n_233, n_234, n_235, n_236, n_237, n_238;
  wire n_239, n_240, n_241, n_242, n_243, n_244, n_245, n_246;
  wire n_247, n_248, n_249, n_250, n_251, n_252, n_253, n_254;
  wire n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_262;
  wire n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270;
  wire n_271, n_272, n_273, n_274, n_275, n_276, n_277, n_278;
  wire n_279, n_280, n_281, n_282, n_283, n_284, n_285, n_286;
  wire n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_294;
  wire n_295, n_296, n_297, n_298, n_299, n_300, n_301, n_302;
  wire n_303, n_304, n_305, n_306, n_307, n_308, n_309, n_310;
  wire n_311, n_312, n_313, n_314, n_315, n_316, n_317, n_318;
  wire n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326;
  wire n_327, n_328, n_329, n_330, n_331, n_332, n_333, n_334;
  wire n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342;
  wire n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350;
  wire n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358;
  wire n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366;
  wire n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374;
  wire n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382;
  wire n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390;
  wire n_391, n_392, n_393, n_394, n_395, n_396, n_397, n_398;
  wire n_399, n_400, n_401, n_402, n_403, n_404, n_405, n_406;
  wire n_407, n_408, n_409, n_410, n_411, n_412, n_413, n_414;
  wire n_415, n_416, n_417, n_418, n_419, n_420, n_421, n_422;
  wire n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430;
  wire n_431, n_432, n_433, n_434, n_435, n_436, n_440;
  nand g1 (n_167, A[0], B[0]);
  nand g2 (n_168, A[0], CI);
  nand g3 (n_169, B[0], CI);
  nand g4 (n_171, n_167, n_168, n_169);
  xor g5 (n_170, A[0], B[0]);
  xor g6 (Z[0], CI, n_170);
  nand g7 (n_172, A[1], B[1]);
  nand g8 (n_173, A[1], n_171);
  nand g9 (n_174, B[1], n_171);
  nand g10 (n_176, n_172, n_173, n_174);
  xor g11 (n_175, A[1], B[1]);
  xor g12 (Z[1], n_171, n_175);
  nand g13 (n_177, A[2], B[2]);
  nand g14 (n_178, A[2], n_176);
  nand g15 (n_179, B[2], n_176);
  nand g16 (n_181, n_177, n_178, n_179);
  xor g17 (n_180, A[2], B[2]);
  xor g18 (Z[2], n_176, n_180);
  nand g19 (n_182, A[3], B[3]);
  nand g20 (n_183, A[3], n_181);
  nand g21 (n_184, B[3], n_181);
  nand g22 (n_186, n_182, n_183, n_184);
  xor g23 (n_185, A[3], B[3]);
  xor g24 (Z[3], n_181, n_185);
  nand g25 (n_187, A[4], B[4]);
  nand g26 (n_188, A[4], n_186);
  nand g27 (n_189, B[4], n_186);
  nand g28 (n_191, n_187, n_188, n_189);
  xor g29 (n_190, A[4], B[4]);
  xor g30 (Z[4], n_186, n_190);
  nand g31 (n_192, A[5], B[5]);
  nand g32 (n_193, A[5], n_191);
  nand g33 (n_194, B[5], n_191);
  nand g34 (n_196, n_192, n_193, n_194);
  xor g35 (n_195, A[5], B[5]);
  xor g36 (Z[5], n_191, n_195);
  nand g37 (n_197, A[6], B[6]);
  nand g38 (n_198, A[6], n_196);
  nand g39 (n_199, B[6], n_196);
  nand g40 (n_201, n_197, n_198, n_199);
  xor g41 (n_200, A[6], B[6]);
  xor g42 (Z[6], n_196, n_200);
  nand g43 (n_202, A[7], B[7]);
  nand g44 (n_203, A[7], n_201);
  nand g45 (n_204, B[7], n_201);
  nand g46 (n_206, n_202, n_203, n_204);
  xor g47 (n_205, A[7], B[7]);
  xor g48 (Z[7], n_201, n_205);
  nand g49 (n_207, A[8], B[8]);
  nand g50 (n_208, A[8], n_206);
  nand g51 (n_209, B[8], n_206);
  nand g52 (n_211, n_207, n_208, n_209);
  xor g53 (n_210, A[8], B[8]);
  xor g54 (Z[8], n_206, n_210);
  nand g55 (n_212, A[9], B[9]);
  nand g56 (n_213, A[9], n_211);
  nand g57 (n_214, B[9], n_211);
  nand g58 (n_216, n_212, n_213, n_214);
  xor g59 (n_215, A[9], B[9]);
  xor g60 (Z[9], n_211, n_215);
  nand g61 (n_217, A[10], B[10]);
  nand g62 (n_218, A[10], n_216);
  nand g63 (n_219, B[10], n_216);
  nand g64 (n_221, n_217, n_218, n_219);
  xor g65 (n_220, A[10], B[10]);
  xor g66 (Z[10], n_216, n_220);
  nand g67 (n_222, A[11], B[11]);
  nand g68 (n_223, A[11], n_221);
  nand g69 (n_224, B[11], n_221);
  nand g70 (n_226, n_222, n_223, n_224);
  xor g71 (n_225, A[11], B[11]);
  xor g72 (Z[11], n_221, n_225);
  nand g73 (n_227, A[12], B[12]);
  nand g74 (n_228, A[12], n_226);
  nand g75 (n_229, B[12], n_226);
  nand g76 (n_231, n_227, n_228, n_229);
  xor g77 (n_230, A[12], B[12]);
  xor g78 (Z[12], n_226, n_230);
  nand g79 (n_232, A[13], B[13]);
  nand g80 (n_233, A[13], n_231);
  nand g81 (n_234, B[13], n_231);
  nand g82 (n_236, n_232, n_233, n_234);
  xor g83 (n_235, A[13], B[13]);
  xor g84 (Z[13], n_231, n_235);
  nand g85 (n_237, A[14], B[14]);
  nand g86 (n_238, A[14], n_236);
  nand g87 (n_239, B[14], n_236);
  nand g88 (n_241, n_237, n_238, n_239);
  xor g89 (n_240, A[14], B[14]);
  xor g90 (Z[14], n_236, n_240);
  nand g91 (n_242, A[15], B[15]);
  nand g92 (n_243, A[15], n_241);
  nand g93 (n_244, B[15], n_241);
  nand g94 (n_246, n_242, n_243, n_244);
  xor g95 (n_245, A[15], B[15]);
  xor g96 (Z[15], n_241, n_245);
  nand g97 (n_247, A[16], B[16]);
  nand g98 (n_248, A[16], n_246);
  nand g99 (n_249, B[16], n_246);
  nand g100 (n_251, n_247, n_248, n_249);
  xor g101 (n_250, A[16], B[16]);
  xor g102 (Z[16], n_246, n_250);
  nand g103 (n_252, A[17], B[17]);
  nand g104 (n_253, A[17], n_251);
  nand g105 (n_254, B[17], n_251);
  nand g106 (n_256, n_252, n_253, n_254);
  xor g107 (n_255, A[17], B[17]);
  xor g108 (Z[17], n_251, n_255);
  nand g109 (n_257, A[18], B[18]);
  nand g110 (n_258, A[18], n_256);
  nand g111 (n_259, B[18], n_256);
  nand g112 (n_261, n_257, n_258, n_259);
  xor g113 (n_260, A[18], B[18]);
  xor g114 (Z[18], n_256, n_260);
  nand g115 (n_262, A[19], B[19]);
  nand g116 (n_263, A[19], n_261);
  nand g117 (n_264, B[19], n_261);
  nand g118 (n_266, n_262, n_263, n_264);
  xor g119 (n_265, A[19], B[19]);
  xor g120 (Z[19], n_261, n_265);
  nand g121 (n_267, A[20], B[20]);
  nand g122 (n_268, A[20], n_266);
  nand g123 (n_269, B[20], n_266);
  nand g124 (n_271, n_267, n_268, n_269);
  xor g125 (n_270, A[20], B[20]);
  xor g126 (Z[20], n_266, n_270);
  nand g127 (n_272, A[21], B[21]);
  nand g128 (n_273, A[21], n_271);
  nand g129 (n_274, B[21], n_271);
  nand g130 (n_276, n_272, n_273, n_274);
  xor g131 (n_275, A[21], B[21]);
  xor g132 (Z[21], n_271, n_275);
  nand g133 (n_277, A[22], B[22]);
  nand g134 (n_278, A[22], n_276);
  nand g135 (n_279, B[22], n_276);
  nand g136 (n_281, n_277, n_278, n_279);
  xor g137 (n_280, A[22], B[22]);
  xor g138 (Z[22], n_276, n_280);
  nand g139 (n_282, A[23], B[23]);
  nand g140 (n_283, A[23], n_281);
  nand g141 (n_284, B[23], n_281);
  nand g142 (n_286, n_282, n_283, n_284);
  xor g143 (n_285, A[23], B[23]);
  xor g144 (Z[23], n_281, n_285);
  nand g145 (n_287, A[24], B[24]);
  nand g146 (n_288, A[24], n_286);
  nand g147 (n_289, B[24], n_286);
  nand g148 (n_291, n_287, n_288, n_289);
  xor g149 (n_290, A[24], B[24]);
  xor g150 (Z[24], n_286, n_290);
  nand g151 (n_292, A[25], B[25]);
  nand g152 (n_293, A[25], n_291);
  nand g153 (n_294, B[25], n_291);
  nand g154 (n_296, n_292, n_293, n_294);
  xor g155 (n_295, A[25], B[25]);
  xor g156 (Z[25], n_291, n_295);
  nand g157 (n_297, A[26], B[26]);
  nand g158 (n_298, A[26], n_296);
  nand g159 (n_299, B[26], n_296);
  nand g160 (n_301, n_297, n_298, n_299);
  xor g161 (n_300, A[26], B[26]);
  xor g162 (Z[26], n_296, n_300);
  nand g163 (n_302, A[27], B[27]);
  nand g164 (n_303, A[27], n_301);
  nand g165 (n_304, B[27], n_301);
  nand g166 (n_306, n_302, n_303, n_304);
  xor g167 (n_305, A[27], B[27]);
  xor g168 (Z[27], n_301, n_305);
  nand g169 (n_307, A[28], B[28]);
  nand g170 (n_308, A[28], n_306);
  nand g171 (n_309, B[28], n_306);
  nand g172 (n_311, n_307, n_308, n_309);
  xor g173 (n_310, A[28], B[28]);
  xor g174 (Z[28], n_306, n_310);
  nand g175 (n_312, A[29], B[29]);
  nand g176 (n_313, A[29], n_311);
  nand g177 (n_314, B[29], n_311);
  nand g178 (n_316, n_312, n_313, n_314);
  xor g179 (n_315, A[29], B[29]);
  xor g180 (Z[29], n_311, n_315);
  nand g181 (n_317, A[30], B[30]);
  nand g182 (n_318, A[30], n_316);
  nand g183 (n_319, B[30], n_316);
  nand g184 (n_321, n_317, n_318, n_319);
  xor g185 (n_320, A[30], B[30]);
  xor g186 (Z[30], n_316, n_320);
  nand g187 (n_322, A[31], B[31]);
  nand g188 (n_323, A[31], n_321);
  nand g189 (n_324, B[31], n_321);
  nand g190 (n_326, n_322, n_323, n_324);
  xor g191 (n_325, A[31], B[31]);
  xor g192 (Z[31], n_321, n_325);
  nand g193 (n_327, A[32], B[32]);
  nand g194 (n_328, A[32], n_326);
  nand g195 (n_329, B[32], n_326);
  nand g196 (n_331, n_327, n_328, n_329);
  xor g197 (n_330, A[32], B[32]);
  xor g198 (Z[32], n_326, n_330);
  nand g199 (n_332, A[33], B[33]);
  nand g200 (n_333, A[33], n_331);
  nand g201 (n_334, B[33], n_331);
  nand g202 (n_336, n_332, n_333, n_334);
  xor g203 (n_335, A[33], B[33]);
  xor g204 (Z[33], n_331, n_335);
  nand g205 (n_337, A[34], B[34]);
  nand g206 (n_338, A[34], n_336);
  nand g207 (n_339, B[34], n_336);
  nand g208 (n_341, n_337, n_338, n_339);
  xor g209 (n_340, A[34], B[34]);
  xor g210 (Z[34], n_336, n_340);
  nand g211 (n_342, A[35], B[35]);
  nand g212 (n_343, A[35], n_341);
  nand g213 (n_344, B[35], n_341);
  nand g214 (n_346, n_342, n_343, n_344);
  xor g215 (n_345, A[35], B[35]);
  xor g216 (Z[35], n_341, n_345);
  nand g217 (n_347, A[36], B[36]);
  nand g218 (n_348, A[36], n_346);
  nand g219 (n_349, B[36], n_346);
  nand g220 (n_351, n_347, n_348, n_349);
  xor g221 (n_350, A[36], B[36]);
  xor g222 (Z[36], n_346, n_350);
  nand g223 (n_352, A[37], B[37]);
  nand g224 (n_353, A[37], n_351);
  nand g225 (n_354, B[37], n_351);
  nand g226 (n_356, n_352, n_353, n_354);
  xor g227 (n_355, A[37], B[37]);
  xor g228 (Z[37], n_351, n_355);
  nand g229 (n_357, A[38], B[38]);
  nand g230 (n_358, A[38], n_356);
  nand g231 (n_359, B[38], n_356);
  nand g232 (n_361, n_357, n_358, n_359);
  xor g233 (n_360, A[38], B[38]);
  xor g234 (Z[38], n_356, n_360);
  nand g235 (n_362, A[39], B[39]);
  nand g236 (n_363, A[39], n_361);
  nand g237 (n_364, B[39], n_361);
  nand g238 (n_366, n_362, n_363, n_364);
  xor g239 (n_365, A[39], B[39]);
  xor g240 (Z[39], n_361, n_365);
  nand g241 (n_367, A[40], B[40]);
  nand g242 (n_368, A[40], n_366);
  nand g243 (n_369, B[40], n_366);
  nand g244 (n_371, n_367, n_368, n_369);
  xor g245 (n_370, A[40], B[40]);
  xor g246 (Z[40], n_366, n_370);
  nand g247 (n_372, A[41], B[41]);
  nand g248 (n_373, A[41], n_371);
  nand g249 (n_374, B[41], n_371);
  nand g250 (n_376, n_372, n_373, n_374);
  xor g251 (n_375, A[41], B[41]);
  xor g252 (Z[41], n_371, n_375);
  nand g253 (n_377, A[42], B[42]);
  nand g254 (n_378, A[42], n_376);
  nand g255 (n_379, B[42], n_376);
  nand g256 (n_381, n_377, n_378, n_379);
  xor g257 (n_380, A[42], B[42]);
  xor g258 (Z[42], n_376, n_380);
  nand g259 (n_382, A[43], B[43]);
  nand g260 (n_383, A[43], n_381);
  nand g261 (n_384, B[43], n_381);
  nand g262 (n_386, n_382, n_383, n_384);
  xor g263 (n_385, A[43], B[43]);
  xor g264 (Z[43], n_381, n_385);
  nand g265 (n_387, A[44], B[44]);
  nand g266 (n_388, A[44], n_386);
  nand g267 (n_389, B[44], n_386);
  nand g268 (n_391, n_387, n_388, n_389);
  xor g269 (n_390, A[44], B[44]);
  xor g270 (Z[44], n_386, n_390);
  nand g271 (n_392, A[45], B[45]);
  nand g272 (n_393, A[45], n_391);
  nand g273 (n_394, B[45], n_391);
  nand g274 (n_396, n_392, n_393, n_394);
  xor g275 (n_395, A[45], B[45]);
  xor g276 (Z[45], n_391, n_395);
  nand g277 (n_397, A[46], B[46]);
  nand g278 (n_398, A[46], n_396);
  nand g279 (n_399, B[46], n_396);
  nand g280 (n_401, n_397, n_398, n_399);
  xor g281 (n_400, A[46], B[46]);
  xor g282 (Z[46], n_396, n_400);
  nand g283 (n_402, A[47], B[47]);
  nand g284 (n_403, A[47], n_401);
  nand g285 (n_404, B[47], n_401);
  nand g286 (n_406, n_402, n_403, n_404);
  xor g287 (n_405, A[47], B[47]);
  xor g288 (Z[47], n_401, n_405);
  nand g289 (n_407, A[48], B[48]);
  nand g290 (n_408, A[48], n_406);
  nand g291 (n_409, B[48], n_406);
  nand g292 (n_411, n_407, n_408, n_409);
  xor g293 (n_410, A[48], B[48]);
  xor g294 (Z[48], n_406, n_410);
  nand g295 (n_412, A[49], B[49]);
  nand g296 (n_413, A[49], n_411);
  nand g297 (n_414, B[49], n_411);
  nand g298 (n_416, n_412, n_413, n_414);
  xor g299 (n_415, A[49], B[49]);
  xor g300 (Z[49], n_411, n_415);
  nand g301 (n_417, A[50], B[50]);
  nand g302 (n_418, A[50], n_416);
  nand g303 (n_419, B[50], n_416);
  nand g304 (n_421, n_417, n_418, n_419);
  xor g305 (n_420, A[50], B[50]);
  xor g306 (Z[50], n_416, n_420);
  nand g307 (n_422, A[51], B[51]);
  nand g308 (n_423, A[51], n_421);
  nand g309 (n_424, B[51], n_421);
  nand g310 (n_426, n_422, n_423, n_424);
  xor g311 (n_425, A[51], B[51]);
  xor g312 (Z[51], n_421, n_425);
  nand g313 (n_427, A[52], B[52]);
  nand g314 (n_428, A[52], n_426);
  nand g315 (n_429, B[52], n_426);
  nand g316 (n_431, n_427, n_428, n_429);
  xor g317 (n_430, A[52], B[52]);
  xor g318 (Z[52], n_426, n_430);
  nand g319 (n_432, A[53], B[53]);
  nand g320 (n_433, A[53], n_431);
  nand g321 (n_434, B[53], n_431);
  nand g322 (n_436, n_432, n_433, n_434);
  xor g323 (n_435, A[53], B[53]);
  xor g324 (Z[53], n_431, n_435);
  xor g329 (n_440, A[54], B[54]);
  xor g330 (Z[54], n_436, n_440);
endmodule

module add_unsigned_carry_2520_GENERIC(A, B, CI, Z);
  input [54:0] A, B;
  input CI;
  output [54:0] Z;
  wire [54:0] A, B;
  wire CI;
  wire [54:0] Z;
  add_unsigned_carry_2520_GENERIC_REAL g1(.A (A), .B (B), .CI (CI), .Z
       (Z));
endmodule

module add_unsigned_carry_2532_GENERIC_REAL(A, B, CI, Z);
// synthesis_equation add_unsigned_carry
  input [65:0] A, B;
  input CI;
  output [65:0] Z;
  wire [65:0] A, B;
  wire CI;
  wire [65:0] Z;
  wire n_200, n_201, n_202, n_203, n_204, n_205, n_206, n_207;
  wire n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_215;
  wire n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223;
  wire n_224, n_225, n_226, n_227, n_228, n_229, n_230, n_231;
  wire n_232, n_233, n_234, n_235, n_236, n_237, n_238, n_239;
  wire n_240, n_241, n_242, n_243, n_244, n_245, n_246, n_247;
  wire n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255;
  wire n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263;
  wire n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_271;
  wire n_272, n_273, n_274, n_275, n_276, n_277, n_278, n_279;
  wire n_280, n_281, n_282, n_283, n_284, n_285, n_286, n_287;
  wire n_288, n_289, n_290, n_291, n_292, n_293, n_294, n_295;
  wire n_296, n_297, n_298, n_299, n_300, n_301, n_302, n_303;
  wire n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_311;
  wire n_312, n_313, n_314, n_315, n_316, n_317, n_318, n_319;
  wire n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327;
  wire n_328, n_329, n_330, n_331, n_332, n_333, n_334, n_335;
  wire n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343;
  wire n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351;
  wire n_352, n_353, n_354, n_355, n_356, n_357, n_358, n_359;
  wire n_360, n_361, n_362, n_363, n_364, n_365, n_366, n_367;
  wire n_368, n_369, n_370, n_371, n_372, n_373, n_374, n_375;
  wire n_376, n_377, n_378, n_379, n_380, n_381, n_382, n_383;
  wire n_384, n_385, n_386, n_387, n_388, n_389, n_390, n_391;
  wire n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399;
  wire n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407;
  wire n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415;
  wire n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423;
  wire n_424, n_425, n_426, n_427, n_428, n_429, n_430, n_431;
  wire n_432, n_433, n_434, n_435, n_436, n_437, n_438, n_439;
  wire n_440, n_441, n_442, n_443, n_444, n_445, n_446, n_447;
  wire n_448, n_449, n_450, n_451, n_452, n_453, n_454, n_455;
  wire n_456, n_457, n_458, n_459, n_460, n_461, n_462, n_463;
  wire n_464, n_465, n_466, n_467, n_468, n_469, n_470, n_471;
  wire n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479;
  wire n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487;
  wire n_488, n_489, n_490, n_491, n_492, n_493, n_494, n_495;
  wire n_496, n_497, n_498, n_499, n_500, n_501, n_502, n_503;
  wire n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511;
  wire n_512, n_513, n_514, n_515, n_516, n_517, n_518, n_519;
  wire n_520, n_521, n_522, n_523, n_524, n_528;
  nand g1 (n_200, A[0], B[0]);
  nand g2 (n_201, A[0], CI);
  nand g3 (n_202, B[0], CI);
  nand g4 (n_204, n_200, n_201, n_202);
  xor g5 (n_203, A[0], B[0]);
  xor g6 (Z[0], CI, n_203);
  nand g7 (n_205, A[1], B[1]);
  nand g8 (n_206, A[1], n_204);
  nand g9 (n_207, B[1], n_204);
  nand g10 (n_209, n_205, n_206, n_207);
  xor g11 (n_208, A[1], B[1]);
  xor g12 (Z[1], n_204, n_208);
  nand g13 (n_210, A[2], B[2]);
  nand g14 (n_211, A[2], n_209);
  nand g15 (n_212, B[2], n_209);
  nand g16 (n_214, n_210, n_211, n_212);
  xor g17 (n_213, A[2], B[2]);
  xor g18 (Z[2], n_209, n_213);
  nand g19 (n_215, A[3], B[3]);
  nand g20 (n_216, A[3], n_214);
  nand g21 (n_217, B[3], n_214);
  nand g22 (n_219, n_215, n_216, n_217);
  xor g23 (n_218, A[3], B[3]);
  xor g24 (Z[3], n_214, n_218);
  nand g25 (n_220, A[4], B[4]);
  nand g26 (n_221, A[4], n_219);
  nand g27 (n_222, B[4], n_219);
  nand g28 (n_224, n_220, n_221, n_222);
  xor g29 (n_223, A[4], B[4]);
  xor g30 (Z[4], n_219, n_223);
  nand g31 (n_225, A[5], B[5]);
  nand g32 (n_226, A[5], n_224);
  nand g33 (n_227, B[5], n_224);
  nand g34 (n_229, n_225, n_226, n_227);
  xor g35 (n_228, A[5], B[5]);
  xor g36 (Z[5], n_224, n_228);
  nand g37 (n_230, A[6], B[6]);
  nand g38 (n_231, A[6], n_229);
  nand g39 (n_232, B[6], n_229);
  nand g40 (n_234, n_230, n_231, n_232);
  xor g41 (n_233, A[6], B[6]);
  xor g42 (Z[6], n_229, n_233);
  nand g43 (n_235, A[7], B[7]);
  nand g44 (n_236, A[7], n_234);
  nand g45 (n_237, B[7], n_234);
  nand g46 (n_239, n_235, n_236, n_237);
  xor g47 (n_238, A[7], B[7]);
  xor g48 (Z[7], n_234, n_238);
  nand g49 (n_240, A[8], B[8]);
  nand g50 (n_241, A[8], n_239);
  nand g51 (n_242, B[8], n_239);
  nand g52 (n_244, n_240, n_241, n_242);
  xor g53 (n_243, A[8], B[8]);
  xor g54 (Z[8], n_239, n_243);
  nand g55 (n_245, A[9], B[9]);
  nand g56 (n_246, A[9], n_244);
  nand g57 (n_247, B[9], n_244);
  nand g58 (n_249, n_245, n_246, n_247);
  xor g59 (n_248, A[9], B[9]);
  xor g60 (Z[9], n_244, n_248);
  nand g61 (n_250, A[10], B[10]);
  nand g62 (n_251, A[10], n_249);
  nand g63 (n_252, B[10], n_249);
  nand g64 (n_254, n_250, n_251, n_252);
  xor g65 (n_253, A[10], B[10]);
  xor g66 (Z[10], n_249, n_253);
  nand g67 (n_255, A[11], B[11]);
  nand g68 (n_256, A[11], n_254);
  nand g69 (n_257, B[11], n_254);
  nand g70 (n_259, n_255, n_256, n_257);
  xor g71 (n_258, A[11], B[11]);
  xor g72 (Z[11], n_254, n_258);
  nand g73 (n_260, A[12], B[12]);
  nand g74 (n_261, A[12], n_259);
  nand g75 (n_262, B[12], n_259);
  nand g76 (n_264, n_260, n_261, n_262);
  xor g77 (n_263, A[12], B[12]);
  xor g78 (Z[12], n_259, n_263);
  nand g79 (n_265, A[13], B[13]);
  nand g80 (n_266, A[13], n_264);
  nand g81 (n_267, B[13], n_264);
  nand g82 (n_269, n_265, n_266, n_267);
  xor g83 (n_268, A[13], B[13]);
  xor g84 (Z[13], n_264, n_268);
  nand g85 (n_270, A[14], B[14]);
  nand g86 (n_271, A[14], n_269);
  nand g87 (n_272, B[14], n_269);
  nand g88 (n_274, n_270, n_271, n_272);
  xor g89 (n_273, A[14], B[14]);
  xor g90 (Z[14], n_269, n_273);
  nand g91 (n_275, A[15], B[15]);
  nand g92 (n_276, A[15], n_274);
  nand g93 (n_277, B[15], n_274);
  nand g94 (n_279, n_275, n_276, n_277);
  xor g95 (n_278, A[15], B[15]);
  xor g96 (Z[15], n_274, n_278);
  nand g97 (n_280, A[16], B[16]);
  nand g98 (n_281, A[16], n_279);
  nand g99 (n_282, B[16], n_279);
  nand g100 (n_284, n_280, n_281, n_282);
  xor g101 (n_283, A[16], B[16]);
  xor g102 (Z[16], n_279, n_283);
  nand g103 (n_285, A[17], B[17]);
  nand g104 (n_286, A[17], n_284);
  nand g105 (n_287, B[17], n_284);
  nand g106 (n_289, n_285, n_286, n_287);
  xor g107 (n_288, A[17], B[17]);
  xor g108 (Z[17], n_284, n_288);
  nand g109 (n_290, A[18], B[18]);
  nand g110 (n_291, A[18], n_289);
  nand g111 (n_292, B[18], n_289);
  nand g112 (n_294, n_290, n_291, n_292);
  xor g113 (n_293, A[18], B[18]);
  xor g114 (Z[18], n_289, n_293);
  nand g115 (n_295, A[19], B[19]);
  nand g116 (n_296, A[19], n_294);
  nand g117 (n_297, B[19], n_294);
  nand g118 (n_299, n_295, n_296, n_297);
  xor g119 (n_298, A[19], B[19]);
  xor g120 (Z[19], n_294, n_298);
  nand g121 (n_300, A[20], B[20]);
  nand g122 (n_301, A[20], n_299);
  nand g123 (n_302, B[20], n_299);
  nand g124 (n_304, n_300, n_301, n_302);
  xor g125 (n_303, A[20], B[20]);
  xor g126 (Z[20], n_299, n_303);
  nand g127 (n_305, A[21], B[21]);
  nand g128 (n_306, A[21], n_304);
  nand g129 (n_307, B[21], n_304);
  nand g130 (n_309, n_305, n_306, n_307);
  xor g131 (n_308, A[21], B[21]);
  xor g132 (Z[21], n_304, n_308);
  nand g133 (n_310, A[22], B[22]);
  nand g134 (n_311, A[22], n_309);
  nand g135 (n_312, B[22], n_309);
  nand g136 (n_314, n_310, n_311, n_312);
  xor g137 (n_313, A[22], B[22]);
  xor g138 (Z[22], n_309, n_313);
  nand g139 (n_315, A[23], B[23]);
  nand g140 (n_316, A[23], n_314);
  nand g141 (n_317, B[23], n_314);
  nand g142 (n_319, n_315, n_316, n_317);
  xor g143 (n_318, A[23], B[23]);
  xor g144 (Z[23], n_314, n_318);
  nand g145 (n_320, A[24], B[24]);
  nand g146 (n_321, A[24], n_319);
  nand g147 (n_322, B[24], n_319);
  nand g148 (n_324, n_320, n_321, n_322);
  xor g149 (n_323, A[24], B[24]);
  xor g150 (Z[24], n_319, n_323);
  nand g151 (n_325, A[25], B[25]);
  nand g152 (n_326, A[25], n_324);
  nand g153 (n_327, B[25], n_324);
  nand g154 (n_329, n_325, n_326, n_327);
  xor g155 (n_328, A[25], B[25]);
  xor g156 (Z[25], n_324, n_328);
  nand g157 (n_330, A[26], B[26]);
  nand g158 (n_331, A[26], n_329);
  nand g159 (n_332, B[26], n_329);
  nand g160 (n_334, n_330, n_331, n_332);
  xor g161 (n_333, A[26], B[26]);
  xor g162 (Z[26], n_329, n_333);
  nand g163 (n_335, A[27], B[27]);
  nand g164 (n_336, A[27], n_334);
  nand g165 (n_337, B[27], n_334);
  nand g166 (n_339, n_335, n_336, n_337);
  xor g167 (n_338, A[27], B[27]);
  xor g168 (Z[27], n_334, n_338);
  nand g169 (n_340, A[28], B[28]);
  nand g170 (n_341, A[28], n_339);
  nand g171 (n_342, B[28], n_339);
  nand g172 (n_344, n_340, n_341, n_342);
  xor g173 (n_343, A[28], B[28]);
  xor g174 (Z[28], n_339, n_343);
  nand g175 (n_345, A[29], B[29]);
  nand g176 (n_346, A[29], n_344);
  nand g177 (n_347, B[29], n_344);
  nand g178 (n_349, n_345, n_346, n_347);
  xor g179 (n_348, A[29], B[29]);
  xor g180 (Z[29], n_344, n_348);
  nand g181 (n_350, A[30], B[30]);
  nand g182 (n_351, A[30], n_349);
  nand g183 (n_352, B[30], n_349);
  nand g184 (n_354, n_350, n_351, n_352);
  xor g185 (n_353, A[30], B[30]);
  xor g186 (Z[30], n_349, n_353);
  nand g187 (n_355, A[31], B[31]);
  nand g188 (n_356, A[31], n_354);
  nand g189 (n_357, B[31], n_354);
  nand g190 (n_359, n_355, n_356, n_357);
  xor g191 (n_358, A[31], B[31]);
  xor g192 (Z[31], n_354, n_358);
  nand g193 (n_360, A[32], B[32]);
  nand g194 (n_361, A[32], n_359);
  nand g195 (n_362, B[32], n_359);
  nand g196 (n_364, n_360, n_361, n_362);
  xor g197 (n_363, A[32], B[32]);
  xor g198 (Z[32], n_359, n_363);
  nand g199 (n_365, A[33], B[33]);
  nand g200 (n_366, A[33], n_364);
  nand g201 (n_367, B[33], n_364);
  nand g202 (n_369, n_365, n_366, n_367);
  xor g203 (n_368, A[33], B[33]);
  xor g204 (Z[33], n_364, n_368);
  nand g205 (n_370, A[34], B[34]);
  nand g206 (n_371, A[34], n_369);
  nand g207 (n_372, B[34], n_369);
  nand g208 (n_374, n_370, n_371, n_372);
  xor g209 (n_373, A[34], B[34]);
  xor g210 (Z[34], n_369, n_373);
  nand g211 (n_375, A[35], B[35]);
  nand g212 (n_376, A[35], n_374);
  nand g213 (n_377, B[35], n_374);
  nand g214 (n_379, n_375, n_376, n_377);
  xor g215 (n_378, A[35], B[35]);
  xor g216 (Z[35], n_374, n_378);
  nand g217 (n_380, A[36], B[36]);
  nand g218 (n_381, A[36], n_379);
  nand g219 (n_382, B[36], n_379);
  nand g220 (n_384, n_380, n_381, n_382);
  xor g221 (n_383, A[36], B[36]);
  xor g222 (Z[36], n_379, n_383);
  nand g223 (n_385, A[37], B[37]);
  nand g224 (n_386, A[37], n_384);
  nand g225 (n_387, B[37], n_384);
  nand g226 (n_389, n_385, n_386, n_387);
  xor g227 (n_388, A[37], B[37]);
  xor g228 (Z[37], n_384, n_388);
  nand g229 (n_390, A[38], B[38]);
  nand g230 (n_391, A[38], n_389);
  nand g231 (n_392, B[38], n_389);
  nand g232 (n_394, n_390, n_391, n_392);
  xor g233 (n_393, A[38], B[38]);
  xor g234 (Z[38], n_389, n_393);
  nand g235 (n_395, A[39], B[39]);
  nand g236 (n_396, A[39], n_394);
  nand g237 (n_397, B[39], n_394);
  nand g238 (n_399, n_395, n_396, n_397);
  xor g239 (n_398, A[39], B[39]);
  xor g240 (Z[39], n_394, n_398);
  nand g241 (n_400, A[40], B[40]);
  nand g242 (n_401, A[40], n_399);
  nand g243 (n_402, B[40], n_399);
  nand g244 (n_404, n_400, n_401, n_402);
  xor g245 (n_403, A[40], B[40]);
  xor g246 (Z[40], n_399, n_403);
  nand g247 (n_405, A[41], B[41]);
  nand g248 (n_406, A[41], n_404);
  nand g249 (n_407, B[41], n_404);
  nand g250 (n_409, n_405, n_406, n_407);
  xor g251 (n_408, A[41], B[41]);
  xor g252 (Z[41], n_404, n_408);
  nand g253 (n_410, A[42], B[42]);
  nand g254 (n_411, A[42], n_409);
  nand g255 (n_412, B[42], n_409);
  nand g256 (n_414, n_410, n_411, n_412);
  xor g257 (n_413, A[42], B[42]);
  xor g258 (Z[42], n_409, n_413);
  nand g259 (n_415, A[43], B[43]);
  nand g260 (n_416, A[43], n_414);
  nand g261 (n_417, B[43], n_414);
  nand g262 (n_419, n_415, n_416, n_417);
  xor g263 (n_418, A[43], B[43]);
  xor g264 (Z[43], n_414, n_418);
  nand g265 (n_420, A[44], B[44]);
  nand g266 (n_421, A[44], n_419);
  nand g267 (n_422, B[44], n_419);
  nand g268 (n_424, n_420, n_421, n_422);
  xor g269 (n_423, A[44], B[44]);
  xor g270 (Z[44], n_419, n_423);
  nand g271 (n_425, A[45], B[45]);
  nand g272 (n_426, A[45], n_424);
  nand g273 (n_427, B[45], n_424);
  nand g274 (n_429, n_425, n_426, n_427);
  xor g275 (n_428, A[45], B[45]);
  xor g276 (Z[45], n_424, n_428);
  nand g277 (n_430, A[46], B[46]);
  nand g278 (n_431, A[46], n_429);
  nand g279 (n_432, B[46], n_429);
  nand g280 (n_434, n_430, n_431, n_432);
  xor g281 (n_433, A[46], B[46]);
  xor g282 (Z[46], n_429, n_433);
  nand g283 (n_435, A[47], B[47]);
  nand g284 (n_436, A[47], n_434);
  nand g285 (n_437, B[47], n_434);
  nand g286 (n_439, n_435, n_436, n_437);
  xor g287 (n_438, A[47], B[47]);
  xor g288 (Z[47], n_434, n_438);
  nand g289 (n_440, A[48], B[48]);
  nand g290 (n_441, A[48], n_439);
  nand g291 (n_442, B[48], n_439);
  nand g292 (n_444, n_440, n_441, n_442);
  xor g293 (n_443, A[48], B[48]);
  xor g294 (Z[48], n_439, n_443);
  nand g295 (n_445, A[49], B[49]);
  nand g296 (n_446, A[49], n_444);
  nand g297 (n_447, B[49], n_444);
  nand g298 (n_449, n_445, n_446, n_447);
  xor g299 (n_448, A[49], B[49]);
  xor g300 (Z[49], n_444, n_448);
  nand g301 (n_450, A[50], B[50]);
  nand g302 (n_451, A[50], n_449);
  nand g303 (n_452, B[50], n_449);
  nand g304 (n_454, n_450, n_451, n_452);
  xor g305 (n_453, A[50], B[50]);
  xor g306 (Z[50], n_449, n_453);
  nand g307 (n_455, A[51], B[51]);
  nand g308 (n_456, A[51], n_454);
  nand g309 (n_457, B[51], n_454);
  nand g310 (n_459, n_455, n_456, n_457);
  xor g311 (n_458, A[51], B[51]);
  xor g312 (Z[51], n_454, n_458);
  nand g313 (n_460, A[52], B[52]);
  nand g314 (n_461, A[52], n_459);
  nand g315 (n_462, B[52], n_459);
  nand g316 (n_464, n_460, n_461, n_462);
  xor g317 (n_463, A[52], B[52]);
  xor g318 (Z[52], n_459, n_463);
  nand g319 (n_465, A[53], B[53]);
  nand g320 (n_466, A[53], n_464);
  nand g321 (n_467, B[53], n_464);
  nand g322 (n_469, n_465, n_466, n_467);
  xor g323 (n_468, A[53], B[53]);
  xor g324 (Z[53], n_464, n_468);
  nand g325 (n_470, A[54], B[54]);
  nand g326 (n_471, A[54], n_469);
  nand g327 (n_472, B[54], n_469);
  nand g328 (n_474, n_470, n_471, n_472);
  xor g329 (n_473, A[54], B[54]);
  xor g330 (Z[54], n_469, n_473);
  nand g331 (n_475, A[55], B[55]);
  nand g332 (n_476, A[55], n_474);
  nand g333 (n_477, B[55], n_474);
  nand g334 (n_479, n_475, n_476, n_477);
  xor g335 (n_478, A[55], B[55]);
  xor g336 (Z[55], n_474, n_478);
  nand g337 (n_480, A[56], B[56]);
  nand g338 (n_481, A[56], n_479);
  nand g339 (n_482, B[56], n_479);
  nand g340 (n_484, n_480, n_481, n_482);
  xor g341 (n_483, A[56], B[56]);
  xor g342 (Z[56], n_479, n_483);
  nand g343 (n_485, A[57], B[57]);
  nand g344 (n_486, A[57], n_484);
  nand g345 (n_487, B[57], n_484);
  nand g346 (n_489, n_485, n_486, n_487);
  xor g347 (n_488, A[57], B[57]);
  xor g348 (Z[57], n_484, n_488);
  nand g349 (n_490, A[58], B[58]);
  nand g350 (n_491, A[58], n_489);
  nand g351 (n_492, B[58], n_489);
  nand g352 (n_494, n_490, n_491, n_492);
  xor g353 (n_493, A[58], B[58]);
  xor g354 (Z[58], n_489, n_493);
  nand g355 (n_495, A[59], B[59]);
  nand g356 (n_496, A[59], n_494);
  nand g357 (n_497, B[59], n_494);
  nand g358 (n_499, n_495, n_496, n_497);
  xor g359 (n_498, A[59], B[59]);
  xor g360 (Z[59], n_494, n_498);
  nand g361 (n_500, A[60], B[60]);
  nand g362 (n_501, A[60], n_499);
  nand g363 (n_502, B[60], n_499);
  nand g364 (n_504, n_500, n_501, n_502);
  xor g365 (n_503, A[60], B[60]);
  xor g366 (Z[60], n_499, n_503);
  nand g367 (n_505, A[61], B[61]);
  nand g368 (n_506, A[61], n_504);
  nand g369 (n_507, B[61], n_504);
  nand g370 (n_509, n_505, n_506, n_507);
  xor g371 (n_508, A[61], B[61]);
  xor g372 (Z[61], n_504, n_508);
  nand g373 (n_510, A[62], B[62]);
  nand g374 (n_511, A[62], n_509);
  nand g375 (n_512, B[62], n_509);
  nand g376 (n_514, n_510, n_511, n_512);
  xor g377 (n_513, A[62], B[62]);
  xor g378 (Z[62], n_509, n_513);
  nand g379 (n_515, A[63], B[63]);
  nand g380 (n_516, A[63], n_514);
  nand g381 (n_517, B[63], n_514);
  nand g382 (n_519, n_515, n_516, n_517);
  xor g383 (n_518, A[63], B[63]);
  xor g384 (Z[63], n_514, n_518);
  nand g385 (n_520, A[64], B[64]);
  nand g386 (n_521, A[64], n_519);
  nand g387 (n_522, B[64], n_519);
  nand g388 (n_524, n_520, n_521, n_522);
  xor g389 (n_523, A[64], B[64]);
  xor g390 (Z[64], n_519, n_523);
  xor g395 (n_528, A[65], B[65]);
  xor g396 (Z[65], n_524, n_528);
endmodule

module add_unsigned_carry_2532_GENERIC(A, B, CI, Z);
  input [65:0] A, B;
  input CI;
  output [65:0] Z;
  wire [65:0] A, B;
  wire CI;
  wire [65:0] Z;
  add_unsigned_carry_2532_GENERIC_REAL g1(.A (A), .B (B), .CI (CI), .Z
       (Z));
endmodule

