# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2010, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr).
# Local time is now Fri, 3 Dec 2010, 19:32:18.
# Main process id is 27821.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO OAI22_X4
  CLASS core ;
  FOREIGN OAI22_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 3.23 BY 1.4 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.1072 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3367 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 ;
    PORT
      LAYER metal1 ;
        POLYGON 1.91 0.56 2.045 0.56 2.045 0.725 2.67 0.725 2.67 0.56 2.805 0.56 2.805 0.795 1.91 0.795  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.146025 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5187 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 ;
    PORT
      LAYER metal1 ;
        POLYGON 1.645 0.425 3.035 0.425 3.035 0.7 2.91 0.7 2.91 0.495 2.39 0.495 2.39 0.66 2.32 0.66 2.32 0.495 1.715 0.495 1.715 0.66 1.645 0.66  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.1072 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3367 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.56 0.52 0.56 0.52 0.725 1.145 0.725 1.145 0.56 1.28 0.56 1.28 0.795 0.385 0.795  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.14565 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5135 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.15 0.425 1.52 0.425 1.52 0.7 1.39 0.7 1.39 0.495 0.865 0.495 0.865 0.66 0.795 0.66 0.795 0.495 0.22 0.495 0.22 0.66 0.15 0.66  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.406 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5262 LAYER metal1 ;
    ANTENNADIFFAREA 0.5852 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.425 0.865 3.1 0.865 3.1 0.36 1.72 0.36 1.72 0.29 3.17 0.29 3.17 0.935 2.765 0.935 2.765 1.21 2.695 1.21 2.695 0.935 2.005 0.935 2.005 1.21 1.935 1.21 1.935 0.935 1.245 0.935 1.245 1.21 1.175 1.21 1.175 0.935 0.495 0.935 0.495 1.21 0.425 1.21  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.04 0.11 1.04 0.11 1.315 0.795 1.315 0.795 1.04 0.865 1.04 0.865 1.315 1.555 1.315 1.555 1.04 1.625 1.04 1.625 1.315 2.315 1.315 2.315 1.04 2.385 1.04 2.385 1.315 3.075 1.315 3.075 1.04 3.145 1.04 3.145 1.315 3.18 1.315 3.23 1.315 3.23 1.485 3.18 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 3.23 -0.085 3.23 0.085 1.435 0.085 1.435 0.195 1.365 0.195 1.365 0.085 1.055 0.085 1.055 0.195 0.985 0.195 0.985 0.085 0.675 0.085 0.675 0.195 0.605 0.195 0.605 0.085 0.295 0.085 0.295 0.195 0.225 0.195 0.225 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.185 0.115 0.185 0.115 0.26 1.525 0.26 1.525 0.15 3.18 0.15 3.18 0.22 1.595 0.22 1.595 0.33 0.045 0.33  ;
  END
END OAI22_X4

END LIBRARY
#
# End of file
#
