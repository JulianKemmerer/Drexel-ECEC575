# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2011, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on server08.nangate.com for user Giancarlo Franciscatto (gfr).
# Local time is now Thu, 6 Jan 2011, 18:10:28.
# Main process id is 3320.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO AON_BUF_X1
  CLASS core ;
  FOREIGN AON_BUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 1.33 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0378 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1586 LAYER metal1 ;
    ANTENNAGATEAREA 0.011 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.28 0.32 0.28 0.32 0.455 0.615 0.455 0.615 0.525 0.25 0.525  ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.04445 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1833 LAYER metal1 ;
    ANTENNADIFFAREA 0.0242 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.82 0.155 0.89 0.155 0.89 0.79 0.82 0.79  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.755 1.315 1.33 1.315 1.33 1.485 0.755 1.485 0 1.485  ;
    END
  END VDD
  PIN VDDBAK
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.92 0.595 0.92 0.595 0.735 0.73 0.735 0.73 0.92 0.755 0.92 0.94 0.92 0.94 1.12 0.755 1.12 0.385 1.12  ;
    END
  END VDDBAK
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 0.73 0.085 0.73 0.25 0.595 0.25 0.595 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.44 0.595 0.685 0.595 0.685 0.385 0.44 0.385 0.44 0.155 0.51 0.155 0.51 0.315 0.755 0.315 0.755 0.665 0.51 0.665 0.51 0.79 0.44 0.79  ;
  END
END AON_BUF_X1

MACRO AON_BUF_X2
  CLASS core ;
  FOREIGN AON_BUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 1.33 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0133 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0611 LAYER metal1 ;
    ANTENNAGATEAREA 0.011 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.42 0.345 0.42 0.345 0.56 0.25 0.56  ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.0427 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1768 LAYER metal1 ;
    ANTENNADIFFAREA 0.04725 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.82 0.215 0.89 0.215 0.89 0.825 0.82 0.825  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.755 1.315 1.33 1.315 1.33 1.485 0.755 1.485 0 1.485  ;
    END
  END VDD
  PIN VDDBAK
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.375 0.92 0.625 0.92 0.625 0.69 0.695 0.69 0.695 0.92 0.755 0.92 0.925 0.92 0.925 1.12 0.755 1.12 0.375 1.12  ;
    END
  END VDDBAK
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 0.72 0.085 0.72 0.24 0.585 0.24 0.585 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.41 0.155 0.48 0.155 0.48 0.46 0.755 0.46 0.755 0.595 0.48 0.595 0.48 0.79 0.41 0.79  ;
  END
END AON_BUF_X2

MACRO AON_BUF_X4
  CLASS core ;
  FOREIGN AON_BUF_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 1.52 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0343 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1417 LAYER metal1 ;
    ANTENNAGATEAREA 0.011 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.42 0.335 0.42 0.335 0.49 0.655 0.49 0.655 0.56 0.25 0.56  ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.06125 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.208 LAYER metal1 ;
    ANTENNADIFFAREA 0.063 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.865 0.215 0.935 0.215 0.935 0.42 1.08 0.42 1.08 0.56 0.935 0.56 0.935 0.8 0.865 0.8  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.8 1.315 1.52 1.315 1.52 1.485 0.8 1.485 0 1.485  ;
    END
  END VDD
  PIN VDDBAK
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.37 0.92 0.675 0.92 0.675 0.81 0.745 0.81 0.745 0.92 0.8 0.92 1.055 0.92 1.055 0.665 1.125 0.665 1.125 1.12 0.8 1.12 0.37 1.12  ;
    END
  END VDDBAK
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.52 -0.085 1.52 0.085 1.125 0.085 1.125 0.28 1.055 0.28 1.055 0.085 0.78 0.085 0.78 0.24 0.645 0.24 0.645 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.44 0.665 0.73 0.665 0.73 0.375 0.47 0.375 0.47 0.155 0.54 0.155 0.54 0.305 0.8 0.305 0.8 0.735 0.44 0.735  ;
  END
END AON_BUF_X4

MACRO AON_INV_X1
  CLASS core ;
  FOREIGN AON_INV_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 1.14 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0168 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0676 LAYER metal1 ;
    ANTENNAGATEAREA 0.011 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.42 0.56 0.42 0.56 0.56 0.44 0.56  ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.04375 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1807 LAYER metal1 ;
    ANTENNADIFFAREA 0.0231 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.17 0.7 0.17 0.7 0.795 0.63 0.795  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN VDDBAK
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4 0.92 0.44 0.92 0.44 0.69 0.51 0.69 0.51 0.92 0.74 0.92 0.74 1.12 0.4 1.12  ;
    END
  END VDDBAK
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.51 0.085 0.51 0.3 0.44 0.3 0.44 0.085 0 0.085  ;
    END
  END VSS
END AON_INV_X1

MACRO AON_INV_X2
  CLASS core ;
  FOREIGN AON_INV_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 1.14 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.01875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.0225 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.28 0.565 0.28 0.565 0.43 0.44 0.43  ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.0434 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1794 LAYER metal1 ;
    ANTENNADIFFAREA 0.04725 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.165 0.7 0.165 0.7 0.785 0.63 0.785  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN VDDBAK
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.395 0.92 0.445 0.92 0.445 0.55 0.515 0.55 0.515 0.92 0.745 0.92 0.745 1.12 0.395 1.12  ;
    END
  END VDDBAK
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.545 0.085 0.545 0.175 0.41 0.175 0.41 0.085 0 0.085  ;
    END
  END VSS
END AON_INV_X2

MACRO AON_INV_X4
  CLASS core ;
  FOREIGN AON_INV_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 1.33 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.019375 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0728 LAYER metal1 ;
    ANTENNAGATEAREA 0.045 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.44 0.28 0.565 0.28 0.565 0.435 0.44 0.435  ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.04375 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1807 LAYER metal1 ;
    ANTENNADIFFAREA 0.06525 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.165 0.7 0.165 0.7 0.79 0.63 0.79  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN VDDBAK
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.38 0.92 0.435 0.92 0.435 0.565 0.505 0.565 0.505 0.92 0.82 0.92 0.82 0.565 0.89 0.565 0.89 0.92 0.95 0.92 0.95 1.12 0.38 1.12  ;
    END
  END VDDBAK
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 0.89 0.085 0.89 0.21 0.82 0.21 0.82 0.085 0.505 0.085 0.505 0.21 0.435 0.21 0.435 0.085 0 0.085  ;
    END
  END VSS
END AON_INV_X4

MACRO HEADER_OE_X1
  CLASS core ;
  FOREIGN HEADER_OE_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 0.95 BY 1.4 ;
  PIN SLEEP
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0595 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1469 LAYER metal1 ;
    ANTENNAGATEAREA 0.018 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.15 0.56 0.575 0.56 0.575 0.7 0.15 0.7  ;
    END
  END SLEEP
  PIN SLEEPOUT
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.0595 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2392 LAYER metal1 ;
    ANTENNADIFFAREA 0.027 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.82 0.18 0.89 0.18 0.89 1.03 0.82 1.03  ;
    END
  END SLEEPOUT
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.115 0.115 1.115 0.115 1.315 0.58 1.315 0.58 0.99 0.715 0.99 0.715 1.315 0.75 1.315 0.95 1.315 0.95 1.485 0.75 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.715 0.085 0.715 0.265 0.58 0.265 0.58 0.085 0 0.085  ;
    END
  END VSS
  PIN VVDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.23 0.84 0.32 0.84 0.32 1.19 0.23 1.19  ;
    END
  END VVDD
  OBS
      LAYER metal1 ;
        POLYGON 0.425 0.835 0.68 0.835 0.68 0.45 0.425 0.45 0.425 0.18 0.495 0.18 0.495 0.38 0.75 0.38 0.75 0.905 0.495 0.905 0.495 1.03 0.425 1.03  ;
  END
END HEADER_OE_X1

MACRO HEADER_OE_X2
  CLASS core ;
  FOREIGN HEADER_OE_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 0.95 BY 1.4 ;
  PIN SLEEP
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0567 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1417 LAYER metal1 ;
    ANTENNAGATEAREA 0.02475 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.15 0.56 0.555 0.56 0.555 0.7 0.15 0.7  ;
    END
  END SLEEP
  PIN SLEEPOUT
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.096425 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2886 LAYER metal1 ;
    ANTENNADIFFAREA 0.05175 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.795 0.165 0.89 0.165 0.89 1.18 0.795 1.18  ;
    END
  END SLEEPOUT
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 0.96 0.11 0.96 0.11 1.315 0.595 1.315 0.595 1.1 0.665 1.1 0.665 1.315 0.725 1.315 0.95 1.315 0.95 1.485 0.725 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.665 0.085 0.665 0.285 0.595 0.285 0.595 0.085 0 0.085  ;
    END
  END VSS
  PIN VVDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.23 0.84 0.32 0.84 0.32 1.18 0.23 1.18  ;
    END
  END VVDD
  OBS
      LAYER metal1 ;
        POLYGON 0.41 0.84 0.655 0.84 0.655 0.425 0.41 0.425 0.41 0.165 0.48 0.165 0.48 0.355 0.725 0.355 0.725 0.91 0.48 0.91 0.48 1.175 0.41 1.175  ;
  END
END HEADER_OE_X2

MACRO HEADER_OE_X4
  CLASS core ;
  FOREIGN HEADER_OE_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 0.95 BY 1.4 ;
  PIN SLEEP
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0466 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1742 LAYER metal1 ;
    ANTENNAGATEAREA 0.03825 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.13 0.42 0.13 0.48 0.59 0.48 0.59 0.56 0.06 0.56  ;
    END
  END SLEEP
  PIN SLEEPOUT
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.06885 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2223 LAYER metal1 ;
    ANTENNADIFFAREA 0.1035 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.8 0.25 0.89 0.25 0.89 1.015 0.8 1.015  ;
    END
  END SLEEPOUT
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 0.985 0.115 0.985 0.115 1.315 0.57 1.315 0.57 0.8 0.705 0.8 0.705 1.315 0.73 1.315 0.95 1.315 0.95 1.485 0.73 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.67 0.085 0.67 0.24 0.6 0.24 0.6 0.085 0 0.085  ;
    END
  END VSS
  PIN VVDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.23 0.7 0.32 0.7 0.32 1.03 0.23 1.03  ;
    END
  END VVDD
  OBS
      LAYER metal1 ;
        POLYGON 0.405 0.66 0.66 0.66 0.66 0.395 0.38 0.395 0.38 0.155 0.515 0.155 0.515 0.325 0.73 0.325 0.73 0.73 0.475 0.73 0.475 0.85 0.405 0.85  ;
  END
END HEADER_OE_X4

MACRO HEADER_X1
  CLASS core ;
  FOREIGN HEADER_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 0.38 BY 1.4 ;
  PIN SLEEP
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.025625 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0858 LAYER metal1 ;
    ANTENNAGATEAREA 0.00675 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.185 0.56 0.185 0.765 0.06 0.765  ;
    END
  END SLEEP
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.005 0.11 1.005 0.11 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0 0.085  ;
    END
  END VSS
  PIN VVDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.23 0.84 0.32 0.84 0.32 1.12 0.23 1.12  ;
    END
  END VVDD
END HEADER_X1

MACRO HEADER_X2
  CLASS core ;
  FOREIGN HEADER_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 0.38 BY 1.4 ;
  PIN SLEEP
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.025625 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0858 LAYER metal1 ;
    ANTENNAGATEAREA 0.0135 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.185 0.56 0.185 0.765 0.06 0.765  ;
    END
  END SLEEP
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 0.96 0.11 0.96 0.11 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0 0.085  ;
    END
  END VSS
  PIN VVDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.23 0.84 0.32 0.84 0.32 1.18 0.23 1.18  ;
    END
  END VVDD
END HEADER_X2

MACRO HEADER_X4
  CLASS core ;
  FOREIGN HEADER_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 0.38 BY 1.4 ;
  PIN SLEEP
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.025625 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0858 LAYER metal1 ;
    ANTENNAGATEAREA 0.027 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.28 0.185 0.28 0.185 0.485 0.06 0.485  ;
    END
  END SLEEP
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 0.985 0.11 0.985 0.11 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0 0.085  ;
    END
  END VSS
  PIN VVDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.23 0.56 0.32 0.56 0.32 1.12 0.23 1.12  ;
    END
  END VVDD
END HEADER_X4

MACRO ISO_FENCE0N_X1
  CLASS core ;
  FOREIGN ISO_FENCE0N_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 0.76 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.02 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0741 LAYER metal1 ;
    ANTENNAGATEAREA 0.01925 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.185 0.56 0.185 0.72 0.06 0.72  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0702 LAYER metal1 ;
    ANTENNAGATEAREA 0.01925 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.42 0.38 0.42 0.38 0.56 0.25 0.56  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.0891 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2808 LAYER metal1 ;
    ANTENNADIFFAREA 0.0378 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.61 0.165 0.7 0.165 0.7 1.155 0.61 1.155  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.06 0.11 1.06 0.11 1.315 0.415 1.315 0.415 1.06 0.485 1.06 0.485 1.315 0.54 1.315 0.76 1.315 0.76 1.485 0.54 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.485 0.085 0.485 0.22 0.415 0.22 0.415 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.235 0.845 0.47 0.845 0.47 0.355 0.045 0.355 0.045 0.19 0.115 0.19 0.115 0.285 0.54 0.285 0.54 0.915 0.305 0.915 0.305 1.065 0.235 1.065  ;
  END
END ISO_FENCE0N_X1

MACRO ISO_FENCE0N_X2
  CLASS core ;
  FOREIGN ISO_FENCE0N_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 0.76 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.01925 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.185 0.42 0.185 0.56 0.06 0.56  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0702 LAYER metal1 ;
    ANTENNAGATEAREA 0.01925 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.42 0.38 0.42 0.38 0.56 0.25 0.56  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.07065 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2275 LAYER metal1 ;
    ANTENNADIFFAREA 0.0756 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.61 0.175 0.7 0.175 0.7 0.96 0.61 0.96  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 0.99 0.11 0.99 0.11 1.315 0.415 1.315 0.415 0.99 0.485 0.99 0.485 1.315 0.54 1.315 0.76 1.315 0.76 1.485 0.54 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.485 0.085 0.485 0.22 0.415 0.22 0.415 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.235 0.725 0.47 0.725 0.47 0.355 0.045 0.355 0.045 0.19 0.115 0.19 0.115 0.285 0.54 0.285 0.54 0.795 0.305 0.795 0.305 0.995 0.235 0.995  ;
  END
END ISO_FENCE0N_X2

MACRO ISO_FENCE0N_X4
  CLASS core ;
  FOREIGN ISO_FENCE0N_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 0.95 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.0365 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.185 0.56 0.185 0.7 0.06 0.7  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0217 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0767 LAYER metal1 ;
    ANTENNAGATEAREA 0.0365 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.56 0.405 0.56 0.405 0.7 0.25 0.7  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.0658 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2626 LAYER metal1 ;
    ANTENNADIFFAREA 0.1008 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.15 0.7 0.15 0.7 1.09 0.63 1.09  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.065 1.315 0.065 0.96 0.135 0.96 0.135 1.315 0.44 1.315 0.44 0.96 0.51 0.96 0.51 1.315 0.56 1.315 0.82 1.315 0.82 0.985 0.89 0.985 0.89 1.315 0.95 1.315 0.95 1.485 0.56 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.89 0.085 0.89 0.34 0.82 0.34 0.82 0.085 0.51 0.085 0.51 0.2 0.44 0.2 0.44 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.26 0.825 0.49 0.825 0.49 0.355 0.035 0.355 0.035 0.285 0.56 0.285 0.56 0.895 0.33 0.895 0.33 1.1 0.26 1.1  ;
  END
END ISO_FENCE0N_X4

MACRO ISO_FENCE0_X1
  CLASS core ;
  FOREIGN ISO_FENCE0_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 0.57 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.014 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0624 LAYER metal1 ;
    ANTENNAGATEAREA 0.02025 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.7 0.35 0.7 0.35 0.84 0.25 0.84  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.02025 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.7 0.185 0.7 0.185 0.84 0.06 0.84  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.086725 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3133 LAYER metal1 ;
    ANTENNADIFFAREA 0.04795 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.2 0.32 0.2 0.32 0.49 0.495 0.49 0.495 1.145 0.42 1.145 0.42 0.56 0.235 0.56  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.185 0.11 1.185 0.11 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.485 0.085 0.485 0.255 0.415 0.255 0.415 0.085 0.11 0.085 0.11 0.255 0.04 0.255 0.04 0.085 0 0.085  ;
    END
  END VSS
END ISO_FENCE0_X1

MACRO ISO_FENCE0_X2
  CLASS core ;
  FOREIGN ISO_FENCE0_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 0.57 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0133 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0611 LAYER metal1 ;
    ANTENNAGATEAREA 0.0405 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.26 0.56 0.355 0.56 0.355 0.7 0.26 0.7  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0702 LAYER metal1 ;
    ANTENNAGATEAREA 0.0405 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.19 0.56 0.19 0.7 0.06 0.7  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.08585 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2977 LAYER metal1 ;
    ANTENNADIFFAREA 0.095725 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.23 0.15 0.3 0.15 0.3 0.415 0.51 0.415 0.51 1.015 0.42 1.015 0.42 0.485 0.23 0.485  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.03 0.11 1.03 0.11 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.485 0.085 0.485 0.335 0.415 0.335 0.415 0.085 0.11 0.085 0.11 0.335 0.04 0.335 0.04 0.085 0 0.085  ;
    END
  END VSS
END ISO_FENCE0_X2

MACRO ISO_FENCE0_X4
  CLASS core ;
  FOREIGN ISO_FENCE0_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 0.95 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0204 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0754 LAYER metal1 ;
    ANTENNAGATEAREA 0.081 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.58 0.42 0.7 0.42 0.7 0.59 0.58 0.59  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.12215 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.416 LAYER metal1 ;
    ANTENNAGATEAREA 0.081 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.18 0.56 0.18 0.98 0.735 0.98 0.735 0.65 0.84 0.65 0.84 1.05 0.11 1.05 0.11 0.7 0.06 0.7  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.077325 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2951 LAYER metal1 ;
    ANTENNADIFFAREA 0.1561 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.215 0.285 0.725 0.285 0.725 0.355 0.51 0.355 0.51 0.91 0.435 0.91 0.435 0.355 0.215 0.355  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.055 1.315 0.055 1.18 0.125 1.18 0.125 1.315 0.815 1.315 0.815 1.18 0.885 1.18 0.885 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.88 0.085 0.88 0.36 0.81 0.36 0.81 0.085 0.5 0.085 0.5 0.22 0.43 0.22 0.43 0.085 0.125 0.085 0.125 0.36 0.055 0.36 0.055 0.085 0 0.085  ;
    END
  END VSS
END ISO_FENCE0_X4

MACRO ISO_FENCE1N_X1
  CLASS core ;
  FOREIGN ISO_FENCE1N_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 0.57 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0147 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0637 LAYER metal1 ;
    ANTENNAGATEAREA 0.01925 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.42 0.355 0.42 0.355 0.56 0.25 0.56  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.01925 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.185 0.42 0.185 0.56 0.06 0.56  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.0922 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3224 LAYER metal1 ;
    ANTENNADIFFAREA 0.0476 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.7 0.42 0.7 0.42 0.185 0.51 0.185 0.51 0.77 0.305 0.77 0.305 1.15 0.235 1.15  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.145 0.11 1.145 0.11 1.315 0.415 1.315 0.415 1.145 0.485 1.145 0.485 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.11 0.085 0.11 0.215 0.04 0.215 0.04 0.085 0 0.085  ;
    END
  END VSS
END ISO_FENCE1N_X1

MACRO ISO_FENCE1N_X2
  CLASS core ;
  FOREIGN ISO_FENCE1N_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 0.57 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0147 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0637 LAYER metal1 ;
    ANTENNAGATEAREA 0.03875 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.56 0.355 0.56 0.355 0.7 0.25 0.7  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.03875 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.185 0.56 0.185 0.7 0.06 0.7  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.08895 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3081 LAYER metal1 ;
    ANTENNADIFFAREA 0.0959 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.23 0.77 0.42 0.77 0.42 0.225 0.51 0.225 0.51 0.84 0.3 0.84 0.3 1.13 0.23 1.13  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.015 0.11 1.015 0.11 1.315 0.42 1.315 0.42 1.015 0.49 1.015 0.49 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.11 0.085 0.11 0.355 0.04 0.355 0.04 0.085 0 0.085  ;
    END
  END VSS
END ISO_FENCE1N_X2

MACRO ISO_FENCE1N_X4
  CLASS core ;
  FOREIGN ISO_FENCE1N_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 0.95 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0189 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.0775 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.405 0.7 0.54 0.7 0.54 0.84 0.405 0.84  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.09125 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2886 LAYER metal1 ;
    ANTENNAGATEAREA 0.0775 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.16 0.7 0.32 0.7 0.32 0.905 0.705 0.905 0.705 0.685 0.775 0.685 0.775 0.975 0.16 0.975  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.12985 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5005 LAYER metal1 ;
    ANTENNADIFFAREA 0.1666 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.215 1.04 0.84 1.04 0.84 0.61 0.44 0.61 0.44 0.28 0.51 0.28 0.51 0.54 0.91 0.54 0.91 1.11 0.215 1.11  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.055 1.315 0.055 1.035 0.125 1.035 0.125 1.315 0.43 1.315 0.43 1.175 0.5 1.175 0.5 1.315 0.81 1.315 0.81 1.175 0.88 1.175 0.88 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.88 0.085 0.88 0.41 0.81 0.41 0.81 0.085 0.125 0.085 0.125 0.41 0.055 0.41 0.055 0.085 0 0.085  ;
    END
  END VSS
END ISO_FENCE1N_X4

MACRO ISO_FENCE1_X1
  CLASS core ;
  FOREIGN ISO_FENCE1_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 0.76 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0154 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.065 LAYER metal1 ;
    ANTENNAGATEAREA 0.02025 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.17 0.42 0.17 0.56 0.06 0.56  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0702 LAYER metal1 ;
    ANTENNAGATEAREA 0.02025 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.56 0.38 0.56 0.38 0.7 0.25 0.7  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.0738 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2366 LAYER metal1 ;
    ANTENNADIFFAREA 0.0378 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.61 0.19 0.7 0.19 0.7 1.01 0.61 1.01  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.415 1.315 0.415 1.005 0.485 1.005 0.485 1.315 0.54 1.315 0.76 1.315 0.76 1.485 0.54 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.485 0.085 0.485 0.245 0.415 0.245 0.415 0.085 0.11 0.085 0.11 0.245 0.04 0.245 0.04 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.82 0.47 0.82 0.47 0.42 0.235 0.42 0.235 0.17 0.305 0.17 0.305 0.35 0.54 0.35 0.54 0.89 0.115 0.89 0.115 1.15 0.045 1.15  ;
  END
END ISO_FENCE1_X1

MACRO ISO_FENCE1_X2
  CLASS core ;
  FOREIGN ISO_FENCE1_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 0.76 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.02025 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.185 0.56 0.185 0.7 0.06 0.7  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0217 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0767 LAYER metal1 ;
    ANTENNAGATEAREA 0.02025 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.7 0.405 0.7 0.405 0.84 0.25 0.84  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.056 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2262 LAYER metal1 ;
    ANTENNADIFFAREA 0.0756 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.28 0.7 0.28 0.7 1.08 0.63 1.08  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.44 1.315 0.44 1.145 0.51 1.145 0.51 1.315 0.565 1.315 0.76 1.315 0.76 1.485 0.565 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.51 0.085 0.51 0.325 0.44 0.325 0.44 0.085 0.14 0.085 0.14 0.325 0.07 0.325 0.07 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.035 1.01 0.495 1.01 0.495 0.505 0.26 0.505 0.26 0.225 0.33 0.225 0.33 0.435 0.565 0.435 0.565 1.08 0.035 1.08  ;
  END
END ISO_FENCE1_X2

MACRO ISO_FENCE1_X4
  CLASS core ;
  FOREIGN ISO_FENCE1_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 0.95 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.037 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.185 0.42 0.185 0.56 0.06 0.56  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0702 LAYER metal1 ;
    ANTENNAGATEAREA 0.037 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.42 0.38 0.42 0.38 0.56 0.25 0.56  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.08685 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2743 LAYER metal1 ;
    ANTENNADIFFAREA 0.1008 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.615 0.15 0.705 0.15 0.705 1.115 0.615 1.115  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.415 1.315 0.415 0.995 0.485 0.995 0.485 1.315 0.545 1.315 0.795 1.315 0.795 0.995 0.865 0.995 0.865 1.315 0.95 1.315 0.95 1.485 0.545 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.865 0.085 0.865 0.355 0.795 0.355 0.795 0.085 0.485 0.085 0.485 0.215 0.415 0.215 0.415 0.085 0.11 0.085 0.11 0.355 0.04 0.355 0.04 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.72 0.475 0.72 0.475 0.355 0.2 0.355 0.2 0.285 0.545 0.285 0.545 0.79 0.115 0.79 0.115 1.08 0.045 1.08  ;
  END
END ISO_FENCE1_X4

MACRO LS_HLEN_X1
  CLASS core ;
  FOREIGN LS_HLEN_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.01925 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.56 0.185 0.56 0.185 0.7 0.06 0.7  ;
    END
  END A
  PIN ISOLN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0702 LAYER metal1 ;
    ANTENNAGATEAREA 0.01925 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.42 0.38 0.42 0.38 0.56 0.25 0.56  ;
    END
  END ISOLN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.07515 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2405 LAYER metal1 ;
    ANTENNADIFFAREA 0.0378 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.61 0.165 0.7 0.165 0.7 1 0.61 1  ;
    END
  END Z
  PIN VDDL
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 0.905 0.11 0.905 0.11 1.315 0.415 1.315 0.415 0.905 0.485 0.905 0.485 1.315 0.54 1.315 0.76 1.315 0.76 1.485 0.54 1.485 0 1.485  ;
    END
  END VDDL
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.485 0.085 0.485 0.22 0.415 0.22 0.415 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.235 0.77 0.47 0.77 0.47 0.355 0.045 0.355 0.045 0.19 0.115 0.19 0.115 0.285 0.54 0.285 0.54 0.84 0.305 0.84 0.305 0.95 0.235 0.95  ;
  END
END LS_HLEN_X1

MACRO LS_HLEN_X2
  CLASS core ;
  FOREIGN LS_HLEN_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.01925 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.185 0.42 0.185 0.56 0.06 0.56  ;
    END
  END A
  PIN ISOLN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0702 LAYER metal1 ;
    ANTENNAGATEAREA 0.01925 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.42 0.38 0.42 0.38 0.56 0.25 0.56  ;
    END
  END ISOLN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.07065 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2275 LAYER metal1 ;
    ANTENNADIFFAREA 0.0756 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.61 0.175 0.7 0.175 0.7 0.96 0.61 0.96  ;
    END
  END Z
  PIN VDDL
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 0.99 0.11 0.99 0.11 1.315 0.415 1.315 0.415 0.99 0.485 0.99 0.485 1.315 0.54 1.315 0.76 1.315 0.76 1.485 0.54 1.485 0 1.485  ;
    END
  END VDDL
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.485 0.085 0.485 0.22 0.415 0.22 0.415 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.235 0.63 0.47 0.63 0.47 0.355 0.045 0.355 0.045 0.19 0.115 0.19 0.115 0.285 0.54 0.285 0.54 0.7 0.305 0.7 0.305 0.995 0.235 0.995  ;
  END
END LS_HLEN_X2

MACRO LS_HLEN_X4
  CLASS core ;
  FOREIGN LS_HLEN_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.02125 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0767 LAYER metal1 ;
    ANTENNAGATEAREA 0.0365 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.185 0.42 0.185 0.59 0.06 0.59  ;
    END
  END A
  PIN ISOLN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.02635 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0845 LAYER metal1 ;
    ANTENNAGATEAREA 0.0365 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.42 0.405 0.42 0.405 0.59 0.25 0.59  ;
    END
  END ISOLN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.0539 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2184 LAYER metal1 ;
    ANTENNADIFFAREA 0.1008 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.63 0.15 0.7 0.15 0.7 0.92 0.63 0.92  ;
    END
  END Z
  PIN VDDL
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.065 1.315 0.065 0.79 0.135 0.79 0.135 1.315 0.44 1.315 0.44 0.79 0.51 0.79 0.51 1.315 0.56 1.315 0.82 1.315 0.82 0.815 0.89 0.815 0.89 1.315 0.95 1.315 0.95 1.485 0.56 1.485 0 1.485  ;
    END
  END VDDL
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.89 0.085 0.89 0.34 0.82 0.34 0.82 0.085 0.51 0.085 0.51 0.2 0.44 0.2 0.44 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.26 0.655 0.49 0.655 0.49 0.355 0.035 0.355 0.035 0.285 0.56 0.285 0.56 0.725 0.33 0.725 0.33 0.93 0.26 0.93  ;
  END
END LS_HLEN_X4

MACRO LS_HL_X1
  CLASS core ;
  FOREIGN LS_HL_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0702 LAYER metal1 ;
    ANTENNAGATEAREA 0.018 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.19 0.42 0.19 0.56 0.06 0.56  ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.0621 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2028 LAYER metal1 ;
    ANTENNADIFFAREA 0.0378 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.42 0.165 0.51 0.165 0.51 0.855 0.42 0.855  ;
    END
  END Z
  PIN VDDL
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.225 1.315 0.225 0.78 0.295 0.78 0.295 1.315 0.35 1.315 0.57 1.315 0.57 1.485 0.35 1.485 0 1.485  ;
    END
  END VDDL
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.295 0.085 0.295 0.22 0.225 0.22 0.225 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.625 0.28 0.625 0.28 0.355 0.045 0.355 0.045 0.165 0.115 0.165 0.115 0.285 0.35 0.285 0.35 0.695 0.115 0.695 0.115 0.785 0.045 0.785  ;
  END
END LS_HL_X1

MACRO LS_HL_X2
  CLASS core ;
  FOREIGN LS_HL_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0702 LAYER metal1 ;
    ANTENNAGATEAREA 0.018 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.19 0.42 0.19 0.56 0.06 0.56  ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.07065 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2275 LAYER metal1 ;
    ANTENNADIFFAREA 0.0756 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.42 0.175 0.51 0.175 0.51 0.96 0.42 0.96  ;
    END
  END Z
  PIN VDDL
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.225 1.315 0.225 0.99 0.295 0.99 0.295 1.315 0.35 1.315 0.57 1.315 0.57 1.485 0.35 1.485 0 1.485  ;
    END
  END VDDL
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.295 0.085 0.295 0.22 0.225 0.22 0.225 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.77 0.28 0.77 0.28 0.355 0.045 0.355 0.045 0.165 0.115 0.165 0.115 0.285 0.35 0.285 0.35 0.84 0.115 0.84 0.115 0.995 0.045 0.995  ;
  END
END LS_HL_X2

MACRO LS_HL_X4
  CLASS core ;
  FOREIGN LS_HL_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0702 LAYER metal1 ;
    ANTENNAGATEAREA 0.02 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.19 0.42 0.19 0.56 0.06 0.56  ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.07065 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2275 LAYER metal1 ;
    ANTENNADIFFAREA 0.1008 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.425 0.15 0.515 0.15 0.515 0.935 0.425 0.935  ;
    END
  END Z
  PIN VDDL
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.225 1.315 0.225 0.815 0.295 0.815 0.295 1.315 0.355 1.315 0.605 1.315 0.605 0.815 0.675 0.815 0.675 1.315 0.76 1.315 0.76 1.485 0.355 1.485 0 1.485  ;
    END
  END VDDL
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.675 0.085 0.675 0.36 0.605 0.36 0.605 0.085 0.295 0.085 0.295 0.22 0.225 0.22 0.225 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.68 0.285 0.68 0.285 0.355 0.045 0.355 0.045 0.18 0.115 0.18 0.115 0.285 0.355 0.285 0.355 0.75 0.115 0.75 0.115 1.075 0.045 1.075  ;
  END
END LS_HL_X4

MACRO LS_LHEN_X1
  CLASS core ;
  FOREIGN LS_LHEN_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 2.66 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0308 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1326 LAYER metal1 ;
    ANTENNAGATEAREA 0.014 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.47 0.53 0.47 0.53 0.54 0.32 0.54 0.32 0.7 0.25 0.7  ;
    END
  END A
  PIN ISOLN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.026325 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0858 LAYER metal1 ;
    ANTENNAGATEAREA 0.0275 ;
    PORT
      LAYER metal1 ;
        POLYGON 1.895 0.645 2.03 0.645 2.03 0.84 1.895 0.84  ;
    END
  END ISOLN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.07725 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2873 LAYER metal1 ;
    ANTENNADIFFAREA 0.0336 ;
    PORT
      LAYER metal1 ;
        POLYGON 2.53 0.16 2.605 0.16 2.605 1.19 2.53 1.19  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.695 1.315 1.215 1.315 1.425 1.315 1.425 1.155 1.495 1.155 1.495 1.315 1.955 1.315 1.955 1.05 2.04 1.05 2.04 1.315 2.32 1.315 2.32 1.08 2.455 1.08 2.455 1.315 2.46 1.315 2.66 1.315 2.66 1.485 2.46 1.485 1.215 1.485 0.695 1.485 0 1.485  ;
    END
  END VDD
  PIN VDDL
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.41 0.92 0.55 0.92 0.55 0.74 0.685 0.74 0.685 0.92 0.695 0.92 0.83 0.92 0.83 1.12 0.695 1.12 0.41 1.12  ;
    END
  END VDDL
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.66 -0.085 2.66 0.085 2.42 0.085 2.42 0.295 2.35 0.295 2.35 0.085 1.875 0.085 1.875 0.32 1.805 0.32 1.805 0.085 0.975 0.085 0.975 0.32 0.905 0.32 0.905 0.085 0.62 0.085 0.62 0.27 0.55 0.27 0.55 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.4 0.605 0.625 0.605 0.625 0.405 0.365 0.405 0.365 0.15 0.435 0.15 0.435 0.335 0.695 0.335 0.695 0.675 0.47 0.675 0.47 0.74 0.4 0.74  ;
        POLYGON 0.705 0.165 0.84 0.165 0.84 0.44 1.145 0.44 1.145 0.325 1.215 0.325 1.215 0.51 0.84 0.51 0.84 0.74 0.77 0.74 0.77 0.235 0.705 0.235  ;
        POLYGON 1.245 0.775 1.28 0.775 1.28 0.185 1.35 0.185 1.35 0.775 1.565 0.775 1.565 0.845 1.315 0.845 1.315 1.23 1.245 1.23  ;
        POLYGON 1.38 0.92 1.64 0.92 1.64 0.575 1.435 0.575 1.435 0.185 1.505 0.185 1.505 0.505 2.325 0.505 2.325 0.575 1.71 0.575 1.71 1.23 1.64 1.23 1.64 1.055 1.38 1.055  ;
        POLYGON 2.16 0.935 2.39 0.935 2.39 0.435 1.975 0.435 1.975 0.16 2.045 0.16 2.045 0.365 2.46 0.365 2.46 1.005 2.23 1.005 2.23 1.19 2.16 1.19  ;
  END
END LS_LHEN_X1

MACRO LS_LHEN_X2
  CLASS core ;
  FOREIGN LS_LHEN_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 2.66 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.03325 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1417 LAYER metal1 ;
    ANTENNAGATEAREA 0.011 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.47 0.565 0.47 0.565 0.54 0.32 0.54 0.32 0.7 0.25 0.7  ;
    END
  END A
  PIN ISOLN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0238 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0806 LAYER metal1 ;
    ANTENNAGATEAREA 0.02225 ;
    PORT
      LAYER metal1 ;
        POLYGON 1.86 0.7 2.03 0.7 2.03 0.84 1.86 0.84  ;
    END
  END ISOLN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.06825 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2717 LAYER metal1 ;
    ANTENNADIFFAREA 0.04725 ;
    PORT
      LAYER metal1 ;
        POLYGON 2.53 0.21 2.6 0.21 2.6 1.185 2.53 1.185  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.705 1.315 1.22 1.315 1.435 1.315 1.435 1.155 1.505 1.155 1.505 1.315 1.965 1.315 1.965 1.05 2.035 1.05 2.035 1.315 2.315 1.315 2.315 1.125 2.45 1.125 2.45 1.315 2.46 1.315 2.66 1.315 2.66 1.485 2.46 1.485 1.22 1.485 0.705 1.485 0 1.485  ;
    END
  END VDD
  PIN VDDL
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.415 0.92 0.55 0.92 0.55 0.74 0.685 0.74 0.685 0.92 0.705 0.92 0.83 0.92 0.83 1.12 0.705 1.12 0.415 1.12  ;
    END
  END VDDL
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.66 -0.085 2.66 0.085 2.45 0.085 2.45 0.225 2.315 0.225 2.315 0.085 1.88 0.085 1.88 0.34 1.81 0.34 1.81 0.085 0.98 0.085 0.98 0.335 0.91 0.335 0.91 0.085 0.605 0.085 0.605 0.27 0.535 0.27 0.535 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.395 0.605 0.635 0.605 0.635 0.405 0.345 0.405 0.345 0.15 0.415 0.15 0.415 0.335 0.705 0.335 0.705 0.675 0.465 0.675 0.465 0.795 0.395 0.795  ;
        POLYGON 0.695 0.17 0.845 0.17 0.845 0.54 1.15 0.54 1.15 0.365 1.22 0.365 1.22 0.61 0.845 0.61 0.845 0.795 0.775 0.795 0.775 0.24 0.695 0.24  ;
        POLYGON 1.245 0.77 1.285 0.77 1.285 0.21 1.355 0.21 1.355 0.77 1.575 0.77 1.575 0.84 1.315 0.84 1.315 1.23 1.245 1.23  ;
        POLYGON 1.385 0.92 1.645 0.92 1.645 0.585 1.44 0.585 1.44 0.21 1.51 0.21 1.51 0.515 2.325 0.515 2.325 0.585 1.715 0.585 1.715 1.23 1.645 1.23 1.645 1.055 1.385 1.055  ;
        POLYGON 2.155 0.835 2.39 0.835 2.39 0.44 1.97 0.44 1.97 0.17 2.04 0.17 2.04 0.37 2.46 0.37 2.46 0.905 2.225 0.905 2.225 1.185 2.155 1.185  ;
  END
END LS_LHEN_X2

MACRO LS_LHEN_X4
  CLASS core ;
  FOREIGN LS_LHEN_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 2.66 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0329 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1404 LAYER metal1 ;
    ANTENNAGATEAREA 0.009 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.47 0.56 0.47 0.56 0.54 0.32 0.54 0.32 0.7 0.25 0.7  ;
    END
  END A
  PIN ISOLN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0231 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.0185 ;
    PORT
      LAYER metal1 ;
        POLYGON 1.865 0.7 2.03 0.7 2.03 0.84 1.865 0.84  ;
    END
  END ISOLN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.07175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2847 LAYER metal1 ;
    ANTENNADIFFAREA 0.0987 ;
    PORT
      LAYER metal1 ;
        POLYGON 2.53 0.18 2.6 0.18 2.6 1.205 2.53 1.205  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.695 1.315 1.21 1.315 1.395 1.315 1.395 1.155 1.53 1.155 1.53 1.315 1.96 1.315 1.96 1.1 2.03 1.1 2.03 1.315 2.34 1.315 2.34 1.1 2.41 1.1 2.41 1.315 2.46 1.315 2.66 1.315 2.66 1.485 2.46 1.485 1.21 1.485 0.695 1.485 0 1.485  ;
    END
  END VDD
  PIN VDDL
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.41 0.92 0.555 0.92 0.555 0.74 0.69 0.74 0.69 0.92 0.695 0.92 0.825 0.92 0.825 1.12 0.695 1.12 0.41 1.12  ;
    END
  END VDDL
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.66 -0.085 2.66 0.085 2.44 0.085 2.44 0.245 2.305 0.245 2.305 0.085 1.875 0.085 1.875 0.335 1.805 0.335 1.805 0.085 0.975 0.085 0.975 0.345 0.905 0.345 0.905 0.085 0.605 0.085 0.605 0.27 0.535 0.27 0.535 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.395 0.605 0.625 0.605 0.625 0.405 0.35 0.405 0.35 0.15 0.42 0.15 0.42 0.335 0.695 0.335 0.695 0.675 0.465 0.675 0.465 0.83 0.395 0.83  ;
        POLYGON 0.695 0.175 0.84 0.175 0.84 0.5 1.14 0.5 1.14 0.38 1.21 0.38 1.21 0.57 0.84 0.57 0.84 0.83 0.77 0.83 0.77 0.245 0.695 0.245  ;
        POLYGON 1.235 0.745 1.28 0.745 1.28 0.2 1.35 0.2 1.35 0.745 1.555 0.745 1.555 0.82 1.305 0.82 1.305 1.245 1.235 1.245  ;
        POLYGON 1.375 0.905 1.46 0.905 1.46 0.965 1.62 0.965 1.62 0.54 1.435 0.54 1.435 0.2 1.505 0.2 1.505 0.47 2.32 0.47 2.32 0.54 1.69 0.54 1.69 1.245 1.62 1.245 1.62 1.05 1.375 1.05  ;
        POLYGON 2.15 0.945 2.39 0.945 2.39 0.395 1.96 0.395 1.96 0.155 2.03 0.155 2.03 0.325 2.46 0.325 2.46 1.015 2.22 1.015 2.22 1.225 2.15 1.225  ;
  END
END LS_LHEN_X4

MACRO LS_LH_X1
  CLASS core ;
  FOREIGN LS_LH_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 2.09 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0161 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0663 LAYER metal1 ;
    ANTENNAGATEAREA 0.01125 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.205 0.42 0.32 0.42 0.32 0.56 0.205 0.56  ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.06615 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2639 LAYER metal1 ;
    ANTENNADIFFAREA 0.0336 ;
    PORT
      LAYER metal1 ;
        POLYGON 1.96 0.19 2.03 0.19 2.03 1.135 1.96 1.135  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 1.37 1.315 1.37 1.085 1.44 1.085 1.44 1.315 1.77 1.315 1.77 1.125 1.84 1.125 1.84 1.315 1.89 1.315 2.09 1.315 2.09 1.485 1.89 1.485 0 1.485  ;
    END
  END VDD
  PIN VDDL
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.92 0.59 0.92 0.59 0.675 0.66 0.675 0.66 0.92 0.855 0.92 0.855 1.12 0.385 1.12  ;
    END
  END VDDL
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.09 -0.085 2.09 0.085 1.845 0.085 1.845 0.28 1.77 0.28 1.77 0.085 1.445 0.085 1.445 0.29 1.375 0.29 1.375 0.085 0.66 0.085 0.66 0.28 0.59 0.28 0.59 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.395 0.15 0.465 0.15 0.465 0.35 0.97 0.35 0.97 0.42 0.465 0.42 0.465 0.77 0.395 0.77  ;
        POLYGON 0.74 0.66 1.045 0.66 1.045 0.25 0.755 0.25 0.755 0.18 1.115 0.18 1.115 0.495 1.36 0.495 1.36 0.565 1.115 0.565 1.115 0.73 0.74 0.73  ;
        POLYGON 1.185 0.69 1.43 0.69 1.43 0.425 1.185 0.425 1.185 0.165 1.255 0.165 1.255 0.355 1.5 0.355 1.5 0.76 1.255 0.76 1.255 1.19 1.185 1.19  ;
        POLYGON 1.32 0.84 1.565 0.84 1.565 0.165 1.635 0.165 1.635 0.405 1.89 0.405 1.89 0.54 1.635 0.54 1.635 1.185 1.565 1.185 1.565 0.975 1.32 0.975  ;
  END
END LS_LH_X1

MACRO LS_LH_X2
  CLASS core ;
  FOREIGN LS_LH_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 2.09 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0147 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0637 LAYER metal1 ;
    ANTENNAGATEAREA 0.011 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.215 0.42 0.32 0.42 0.32 0.56 0.215 0.56  ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.07 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2782 LAYER metal1 ;
    ANTENNADIFFAREA 0.04725 ;
    PORT
      LAYER metal1 ;
        POLYGON 1.96 0.215 2.03 0.215 2.03 1.215 1.96 1.215  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 1.41 1.315 1.41 1.085 1.48 1.085 1.48 1.315 1.77 1.315 1.77 0.985 1.84 0.985 1.84 1.315 1.89 1.315 2.09 1.315 2.09 1.485 1.89 1.485 0 1.485  ;
    END
  END VDD
  PIN VDDL
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.92 0.565 0.92 0.565 0.7 0.7 0.7 0.7 0.92 0.88 0.92 0.88 1.12 0.385 1.12  ;
    END
  END VDDL
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.09 -0.085 2.09 0.085 1.84 0.085 1.84 0.28 1.77 0.28 1.77 0.085 1.485 0.085 1.485 0.275 1.415 0.275 1.415 0.085 0.7 0.085 0.7 0.24 0.565 0.24 0.565 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.395 0.15 0.465 0.15 0.465 0.33 1.01 0.33 1.01 0.4 0.465 0.4 0.465 0.77 0.395 0.77  ;
        POLYGON 0.765 0.66 1.08 0.66 1.08 0.25 0.765 0.25 0.765 0.18 1.15 0.18 1.15 0.51 1.395 0.51 1.395 0.58 1.15 0.58 1.15 0.73 0.765 0.73  ;
        POLYGON 1.225 0.695 1.465 0.695 1.465 0.415 1.225 0.415 1.225 0.155 1.295 0.155 1.295 0.345 1.535 0.345 1.535 0.765 1.295 0.765 1.295 1.19 1.225 1.19  ;
        POLYGON 1.36 0.84 1.605 0.84 1.605 0.155 1.675 0.155 1.675 0.495 1.89 0.495 1.89 0.63 1.675 0.63 1.675 1.185 1.605 1.185 1.605 0.975 1.36 0.975  ;
  END
END LS_LH_X2

MACRO LS_LH_X4
  CLASS core ;
  FOREIGN LS_LH_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 2.09 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0168 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0676 LAYER metal1 ;
    ANTENNAGATEAREA 0.011 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2 0.42 0.32 0.42 0.32 0.56 0.2 0.56  ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.05355 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2171 LAYER metal1 ;
    ANTENNADIFFAREA 0.0957 ;
    PORT
      LAYER metal1 ;
        POLYGON 1.96 0.21 2.03 0.21 2.03 0.975 1.96 0.975  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 1.42 1.315 1.42 1.085 1.49 1.085 1.49 1.315 1.765 1.315 1.765 0.985 1.835 0.985 1.835 1.315 1.89 1.315 2.09 1.315 2.09 1.485 1.89 1.485 0 1.485  ;
    END
  END VDD
  PIN VDDL
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.92 0.565 0.92 0.565 0.695 0.7 0.695 0.7 0.92 0.88 0.92 0.88 1.12 0.385 1.12  ;
    END
  END VDDL
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.09 -0.085 2.09 0.085 1.835 0.085 1.835 0.415 1.765 0.415 1.765 0.085 1.495 0.085 1.495 0.275 1.425 0.275 1.425 0.085 0.7 0.085 0.7 0.25 0.565 0.25 0.565 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.395 0.155 0.465 0.155 0.465 0.33 1.01 0.33 1.01 0.4 0.465 0.4 0.465 0.77 0.395 0.77  ;
        POLYGON 0.765 0.665 1.08 0.665 1.08 0.25 0.765 0.25 0.765 0.18 1.15 0.18 1.15 0.5 1.405 0.5 1.405 0.57 1.15 0.57 1.15 0.735 0.765 0.735  ;
        POLYGON 1.235 0.695 1.475 0.695 1.475 0.415 1.235 0.415 1.235 0.155 1.305 0.155 1.305 0.345 1.545 0.345 1.545 0.765 1.305 0.765 1.305 1.19 1.235 1.19  ;
        POLYGON 1.37 0.865 1.615 0.865 1.615 0.155 1.685 0.155 1.685 0.515 1.89 0.515 1.89 0.65 1.685 0.65 1.685 1.185 1.615 1.185 1.615 1.005 1.37 1.005  ;
  END
END LS_LH_X4

END LIBRARY
#
# End of file
#
