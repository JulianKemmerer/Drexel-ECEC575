# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2011, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on server08.nangate.com for user Giancarlo Franciscatto (gfr).
# Local time is now Thu, 6 Jan 2011, 18:10:28.
# Main process id is 3320.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO ISO_FENCE1N_X1
  CLASS core ;
  FOREIGN ISO_FENCE1N_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 0.57 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0147 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0637 LAYER metal1 ;
    ANTENNAGATEAREA 0.01925 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.25 0.42 0.355 0.42 0.355 0.56 0.25 0.56  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.01925 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.06 0.42 0.185 0.42 0.185 0.56 0.06 0.56  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.0922 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3224 LAYER metal1 ;
    ANTENNADIFFAREA 0.0476 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.7 0.42 0.7 0.42 0.185 0.51 0.185 0.51 0.77 0.305 0.77 0.305 1.15 0.235 1.15  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.145 0.11 1.145 0.11 1.315 0.415 1.315 0.415 1.145 0.485 1.145 0.485 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.11 0.085 0.11 0.215 0.04 0.215 0.04 0.085 0 0.085  ;
    END
  END VSS
END ISO_FENCE1N_X1

END LIBRARY
#
# End of file
#
