# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2011, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on server08.nangate.com for user Giancarlo Franciscatto (gfr).
# Local time is now Thu, 6 Jan 2011, 18:10:28.
# Main process id is 3320.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO LS_LH_X4
  CLASS core ;
  FOREIGN LS_LH_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 2.09 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0168 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0676 LAYER metal1 ;
    ANTENNAGATEAREA 0.011 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2 0.42 0.32 0.42 0.32 0.56 0.2 0.56  ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.05355 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2171 LAYER metal1 ;
    ANTENNADIFFAREA 0.0957 ;
    PORT
      LAYER metal1 ;
        POLYGON 1.96 0.21 2.03 0.21 2.03 0.975 1.96 0.975  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 1.42 1.315 1.42 1.085 1.49 1.085 1.49 1.315 1.765 1.315 1.765 0.985 1.835 0.985 1.835 1.315 1.89 1.315 2.09 1.315 2.09 1.485 1.89 1.485 0 1.485  ;
    END
  END VDD
  PIN VDDL
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.92 0.565 0.92 0.565 0.695 0.7 0.695 0.7 0.92 0.88 0.92 0.88 1.12 0.385 1.12  ;
    END
  END VDDL
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.09 -0.085 2.09 0.085 1.835 0.085 1.835 0.415 1.765 0.415 1.765 0.085 1.495 0.085 1.495 0.275 1.425 0.275 1.425 0.085 0.7 0.085 0.7 0.25 0.565 0.25 0.565 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.395 0.155 0.465 0.155 0.465 0.33 1.01 0.33 1.01 0.4 0.465 0.4 0.465 0.77 0.395 0.77  ;
        POLYGON 0.765 0.665 1.08 0.665 1.08 0.25 0.765 0.25 0.765 0.18 1.15 0.18 1.15 0.5 1.405 0.5 1.405 0.57 1.15 0.57 1.15 0.735 0.765 0.735  ;
        POLYGON 1.235 0.695 1.475 0.695 1.475 0.415 1.235 0.415 1.235 0.155 1.305 0.155 1.305 0.345 1.545 0.345 1.545 0.765 1.305 0.765 1.305 1.19 1.235 1.19  ;
        POLYGON 1.37 0.865 1.615 0.865 1.615 0.155 1.685 0.155 1.685 0.515 1.89 0.515 1.89 0.65 1.685 0.65 1.685 1.185 1.615 1.185 1.615 1.005 1.37 1.005  ;
  END
END LS_LH_X4

END LIBRARY
#
# End of file
#
