# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2010, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr).
# Local time is now Fri, 3 Dec 2010, 19:32:18.
# Main process id is 27821.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO SDFFRS_X2
  CLASS core ;
  FOREIGN SDFFRS_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  SIZE 5.89 BY 1.4 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0203 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0741 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 ;
    PORT
      LAYER metal1 ;
        POLYGON 5.495 0.42 5.64 0.42 5.64 0.56 5.495 0.56  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.024025 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0806 LAYER metal1 ;
    ANTENNAGATEAREA 0.075 ;
    PORT
      LAYER metal1 ;
        POLYGON 1.01 0.545 1.165 0.545 1.165 0.7 1.01 0.7  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.07535 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2769 LAYER metal1 ;
    ANTENNAGATEAREA 0.05775 ;
    PORT
      LAYER metal1 ;
        POLYGON 5.135 0.385 5.205 0.385 5.205 0.72 5.57 0.72 5.57 0.675 5.7 0.675 5.7 0.84 5.57 0.84 5.57 0.79 5.135 0.79  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.0203 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0741 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 ;
    PORT
      LAYER metal1 ;
        POLYGON 4.925 0.56 5.07 0.56 5.07 0.7 4.925 0.7  ;
    END
  END SI
  PIN SN
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.014725 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.065 LAYER metal1 ;
    ANTENNAGATEAREA 0.04875 ;
    PORT
      LAYER metal1 ;
        POLYGON 1.365 0.545 1.46 0.545 1.46 0.7 1.365 0.7  ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    ANTENNAPARTIALMETALAREA 0.01155 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0611 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 ;
    PORT
      LAYER metal1 ;
        POLYGON 1.9 0.175 2.065 0.175 2.065 0.245 1.9 0.245  ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2743 LAYER metal1 ;
    ANTENNADIFFAREA 0.1463 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.24 0.15 0.32 0.15 0.32 1.125 0.24 1.125  ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    ANTENNAPARTIALMETALAREA 0.062775 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.156 LAYER metal1 ;
    ANTENNADIFFAREA 0.1463 ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6 0.435 0.735 0.435 0.735 0.9 0.6 0.9  ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.065 1.315 0.065 0.85 0.135 0.85 0.135 1.315 0.41 1.315 0.41 1.1 0.545 1.1 0.545 1.315 0.79 1.315 0.79 1.1 0.925 1.1 0.925 1.315 1.18 1.315 1.18 1.12 1.315 1.12 1.315 1.315 1.64 1.315 1.64 1.115 1.775 1.115 1.775 1.315 2.22 1.315 2.285 1.315 2.285 0.965 2.42 0.965 2.42 1.315 3.04 1.315 3.04 0.985 3.175 0.985 3.175 1.315 3.42 1.315 3.42 0.985 3.555 0.985 3.555 1.315 3.95 1.315 3.95 1.09 4.085 1.09 4.085 1.315 4.24 1.315 4.675 1.315 4.78 1.315 4.78 1.09 4.915 1.09 4.915 1.315 5.295 1.315 5.54 1.315 5.54 1.195 5.675 1.195 5.675 1.315 5.835 1.315 5.89 1.315 5.89 1.485 5.835 1.485 5.295 1.485 4.675 1.485 4.24 1.485 2.22 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 5.89 -0.085 5.89 0.085 5.675 0.085 5.675 0.18 5.54 0.18 5.54 0.085 4.88 0.085 4.88 0.27 4.81 0.27 4.81 0.085 3.895 0.085 3.895 0.285 3.76 0.285 3.76 0.085 3.175 0.085 3.175 0.285 3.04 0.285 3.04 0.085 2.2 0.085 2.2 0.32 2.13 0.32 2.13 0.085 1.835 0.085 1.835 0.285 1.7 0.285 1.7 0.085 0.925 0.085 0.925 0.16 0.79 0.16 0.79 0.085 0.545 0.085 0.545 0.16 0.41 0.16 0.41 0.085 0.135 0.085 0.135 0.41 0.065 0.41 0.065 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.39 0.23 1.305 0.23 1.305 0.3 0.46 0.3 0.46 0.965 1.12 0.965 1.12 1.035 0.39 1.035  ;
        POLYGON 0.94 0.765 1.465 0.765 1.465 0.975 1.91 0.975 1.91 1.16 2.22 1.16 2.22 1.23 1.84 1.23 1.84 1.045 1.395 1.045 1.395 0.835 0.87 0.835 0.87 0.41 1.46 0.41 1.46 0.48 0.94 0.48  ;
        POLYGON 2.13 0.83 2.57 0.83 2.57 1.05 2.5 1.05 2.5 0.9 2.2 0.9 2.2 1.05 2.13 1.05  ;
        POLYGON 1.6 0.84 1.97 0.84 1.97 0.685 2.565 0.685 2.565 0.62 2.635 0.62 2.635 0.755 2.04 0.755 2.04 0.91 1.53 0.91 1.53 0.35 2.04 0.35 2.04 0.42 1.6 0.42  ;
        POLYGON 1.665 0.485 2.7 0.485 2.7 0.2 2.77 0.2 2.77 1.05 2.7 1.05 2.7 0.555 1.735 0.555 1.735 0.68 1.665 0.68  ;
        POLYGON 2.99 0.485 3.455 0.485 3.455 0.32 3.525 0.32 3.525 0.49 4.17 0.49 4.17 0.56 3.06 0.56 3.06 0.765 3.37 0.765 3.37 0.835 2.99 0.835  ;
        POLYGON 3.8 0.955 4.24 0.955 4.24 1.175 4.17 1.175 4.17 1.025 3.87 1.025 3.87 1.175 3.8 1.175  ;
        POLYGON 3.125 0.625 4.405 0.625 4.405 0.285 4.54 0.285 4.54 0.355 4.475 0.355 4.475 0.625 4.51 0.625 4.51 1.09 4.44 1.09 4.44 0.695 3.125 0.695  ;
        POLYGON 3.615 0.765 4.375 0.765 4.375 1.155 4.605 1.155 4.605 0.825 4.575 0.825 4.575 0.69 4.605 0.69 4.605 0.22 4.34 0.22 4.34 0.425 3.61 0.425 3.61 0.22 3.39 0.22 3.39 0.42 2.915 0.42 2.915 1.185 2.555 1.185 2.555 1.115 2.845 1.115 2.845 0.35 3.32 0.35 3.32 0.15 3.68 0.15 3.68 0.355 4.27 0.355 4.27 0.15 4.675 0.15 4.675 1.225 4.305 1.225 4.305 0.835 3.615 0.835  ;
        POLYGON 4.81 0.95 5.295 0.95 5.295 1.02 4.74 1.02 4.74 0.375 4.975 0.375 4.975 0.165 5.295 0.165 5.295 0.235 5.045 0.235 5.045 0.445 4.81 0.445  ;
        POLYGON 5.27 0.565 5.34 0.565 5.34 0.285 5.765 0.285 5.765 0.15 5.835 0.15 5.835 1.09 5.765 1.09 5.765 0.355 5.41 0.355 5.41 0.635 5.27 0.635  ;
  END
END SDFFRS_X2

END LIBRARY
#
# End of file
#
